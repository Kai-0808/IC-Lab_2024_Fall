`define CYCLE_TIME 15.0
`define SEED_NUMBER 19385032
`define PATTERN_NUMBER 10000
`define DEBUG_MODE 1

`include "Usertype.sv"

program automatic PATTERN(input clk, INF.PATTERN inf);

`protected
b^=H8Xd<O)=.>Cd1UgDY1XK_4cf<EMe(1JT-._GOK6d@N)?M@\=>0)E#F<C<#-2#
Nb3f:YU1P2EB3ZZ_CU1Q7JOcQN5=JO05eZ<Hb:7UfFb6PEMAFUa>/]_-6K,gG/B<
^FI1DebU]&b2g,G/ffYUHN=b>]+dE2??eZ5_]9BXc0OeA6g<45M,Q80@W]gCZb_c
4f#49d:aBLdLK+]Gc0:@Q8#]I]gZ^B0L@ZN1ZR&e_NT@:bM&6@^XYcH1MK>+CG&S
HBcgSO576F86[NHbZ-[<f;YH0>W+6=IT)Ua9/3bL??CYb>g=Z0;Da1&R1d>Q\2O1
F3YbB)FZ.f#M^#QW(2/,\YbLJ,4cKLI:MdQ:1dVa#\BAQT01faG8&->#E6@QD,(H
^2GMJ_7U=F=O9D0-P2=R[S(VOXAKWW#Z+R=[YMZ)\JUNdA/Fd6+/6Q^9^U-Weag)
58)>.?+d7g2]/[::6)+C4P^2;[[g#DB@J+^gDR@+#ZF;#ZfL.Z1]>SYL\H+8J8YZ
<-aGVdW-)Z@fB9-c#Q33PCFY7840OdK_Og#e3+1W_OT&4P)25<55-//W&5Qa]g@=
.g#E]<VNXXR4-N;d\51W3:4BHAf\W@&)d&Z8--KX^:X(MOF0X3Z]9H4c(M20:QSW
;#5TL:8LY[YgU)QV7&Be]L_eaS#&3J-=gDM1CUgLAdI,_f4#\H8ML\fR,K[[1/=L
J]\LKLUA@gS<JWDBKIF\KE(+9(#3K[+faR/_0Zc-/>UCH,bc4[>?[?\Ra&8J:ZA.
QD0Sb3ULa1@1cVRUeI1?^JWR8-c<<e^FD,K,WVaaS\[cVNU7^8@^?Ef&^NR&&=gA
V,0bg&34N-B+WgUdg=0MDeEB.&_Qc.H+:/.aZ#(KBCNaVdRP=PHDUPcbRa^3HXQ<
-T_ebO5d6dX93Q2/gP_:+b:WQ->VB,R+3V+D=JO-YM97[(>5WC80YL.S8PYW/O&A
Q?;fAI1YHg&dZE\F&/V])b(^@0B;bM,ZYJbEa[B-gM72-G&_V_QPb8>?MGd?PSY#
-8c8\+2JE4Z40IGb=5F.,KG=0Q71Ce0=McX@;+3AY@HFPg<XQIbIL>?N]C2_F?)_
#/?feQa-E>[YJa>46,/#Vd)&U;@8efNef+R\D.G+=#)QgQX_/\Z(7>gP_F]4BIg,
UZeg\MW+:^4ZY1?A-+5<1@Y2B1fEf)aRF\;G4@3gS3cMU]SKIeG[[d]b.JQ1K_e^
WPF6A[0/a\_gdZJ<@^]3=UE74]2S:,\=][=<&S39;<2KAa/K9;Q:](S>/C5P/d7-
BD&17TUd&Y<b4aH\=4:4#Z86F-\-6YS73.H,3aX)>M:#P_fEF>b>\N2<VD46&J;5
]eLY1G-_Bbc_Lg5NcJC=T.V?aELI=(@X7;3aSGcFO4D519IW<DCNf^C.6L_]fBBA
Xf-;4Z.bY\bRa/91e>-AH?a1E4SC&_W=BLM>:1Y^eP]#e2Ic]A=\)+GA2,<4cV23
S07^QQB&=6XIS<R7W^4NV[f6@W0JC+>\A4@U<;<K0CWH;QW79/A]Af7<90,Vc3MG
IIIbP=O()V8KbV9[aCV;<[<4N9JV9R;=_GMU4]a5ceYF16c[PTc9.cL?dDb<G&U]
IQ4((^2BU&cZg\L#097BLZ+)M]I1ZVD,4Ve)0LJR[ceC;Z9[4.9+:]?GEUg6UA7<
KNF^eWcT8If70M2AbZS0e)Jd8Z^.P==/SCYQEN]Ne.Y9B3<KC(+\TG_/&DAcFJH#
\b#Kf:<2WF[Nba<MQG+0-D-ME+G@bIYY](:[cEC3/O60Qg@Q=eM?T6H>Se:#(3EV
T^HM3(M=BSI(,@+XFHCcCHIM?=1&5+g?GBRf6#0UM_)RAOK[-79@:<PbKO/6Ec#Q
^Y_M<S^-3/]/CB]=#X=FV)(eH:XZL28IBQXJL)A1:<=&CeN8^/F6-aA6:)Gb0[Jf
Jb9cAI/(cAV\B+<EgYb8.Y.-WB29,\GCQYdTA7GD.6T5,6=@1.\:?4<]O58(QIT&
;]<OO:1ME+(V.-\#K4ge,Y./E.<E<f^JcB,F@f548a33LD>7LBRL2_7Z=&+4\W8c
^X=:8aGGO?cD9-CQM[XI)>-dcTBY6FHaH.]9Q0W^YL6[Z<4dQK21+&UF2.88NH1C
2dL7Y1;I?+P[RXGGCeYfD^ZDHEN@NF=1J5#3GaRLBadT-O+1E/Q969ZB:E4M@9Hg
#<&;V/[[)PBfLJY1(]GAF7<8EE;\K?f/#>/bBF.4B#))L)>FK+7Q7/ZKEE+dFbR3
+0_)-CD,Jb,ARM3TX8gBOPSQ>4VNW8@WCcbO>7cT6#\S<gQAZ#]61^0YNY1[@HL(
\5#4DPOc4<@e3H-(M@d3Ae5C<b(TV6&\K#/Oa_08SY/6\94X1B.e\d3LC#aUH\@Y
4c+:eF-,A#=cSQ.#F+_131FRFf=[)=FS2^8_JKQe/a4N-#_W&_^1KDDT:2e3FDRa
#<DCP4+f;L(I]59JJ;S7@Cb7[HBH:8RZ,:(cIKV&WI(<IVNFZC,Z.d@K:VG4^S6B
ATFQ[Z/^=6P/;B;=.;WCZVTS&-;J;K:5W>8=.6[[<S\@,RH6Z]?c++Q7THf57/WK
_;ZI[dda^R?^M#@(9(4_X;Sg).80J:5S#-@_M0-dgCeULW[4[UF.S5R9@7G9]0+c
INWCMR?/d:BeBJB1f]5JdU:0(\E95^A[&QCddB,U6W@WLD=(1D;1=faU[4K-fO_]
eE7?XCQ-B7X@)#0fKOL0fKMQN&d;XGI6F_DSf&,Z.5]R)E^TK,B3TLBAcaeHROUa
8GEE4]89a=e@HK-&5a\.B=g5A<&XB\M+4LK]8EO5O[)L=<:&H][COXaD0adV(>3E
+7+#(53+\#<c4VRdFge]N6/g0aX]&Fg[#Y;KMV=H\+\M9X6(Y#H&H#^;DPX;37/I
B?c<8[H[M2E6a9BW8D.^#COa;I-&.YfK:O+OTG96/(XKUY^A,?9F&@+Gd4&GLVY0
b.FUM<eZV?0Y/@AT^S^F@WJ;;R#HBa=P/:S[+:W,:1#<)bM;eaZV7K];CJb)BSI+
,9A6VW3Y/\\L8&)1Ta93HGBC>^?82/Og-cGTV.S?&];UbEY,7-g/G]HDK6NOLXS+
-+SZ\f(30<g=N(6.X2#U&]DM)Ie044@6e[5<)FU5:==bYa67+E4>F[STYbMV6LL:
:?MNWBW&-765:EV/\MW?8>^<=f&Nf05cS#6MI:4:LOSG,VLLRRO<^I+O1Ff9Nd0c
b-+(=0G:@\/CW^AM33NV]cYc7eO^:U87OG9G=H-cQ7M_<4?T@DO(V-QedQM2F;\@
Hgf73)5./[)BdOE\UA?8PY[IE7GcV)I@L9X;JN4?:,HcO8R]1Y2bJ_GW=&TO&+^[
D533:Z5RC2=/(eF_.X>X#6b[>L_J.BQaB)@O=3Z1AYd3+YZWKVJG+6A6)(XRg4GG
?,UV.bXFSD;Te-4H\8S>(4JeTW]46++156;U;LQ>A?UTeHfgeZ)]b5G3JX;^MQ,6
GQU,^^LDK-UETMT=M[[H.:5-SL.1a8ARX]G^\,g@5EW?81\f]dT8NW._@@IGE6I4
:_=M)a8V?I-PJ9S6_+0=WKL(_1E#JTXFUdYYSbG?T^T?_S0MI3ab&SO0eR8148g0
VUe69f^(E)YA_RMKDS@Pg5^3c/+JD>PKKgR-e_Mb77A?;3Q#_QDZCSJO_fQO?^a8
bJUKNE/OX_=Q[Z?_aWYD(5I;g?/U>;[D&:01=/P\R\g_d;4V]#&U<]9/TAWI<JOA
81KeD7EE:Z^Y?@JP@3+ceOPSD3G<SOD]7BI@FSKfQ=^_9=JM@,X=QOLF0O02:]a?
L/7ER#BFON]-L=PN.TU)7d,]fSb?SC@Oa</)-^T17+L\QFB4/HH.@J5KBB=?I,[C
UYVc+6^M,1fKOS6C=RP@E7<@gbeSFI1I7)F0M#C/]]W/FT\_J.9;,#]eUWN\@)V1
71fW](O+Z.-a&;04QP+6OY477eKCY119+HEBQU_[;ZC8d>^Y[IAKXX]2#;\1WS,f
2S\e+>^?@eU,HJZ#6Z7WDZ[<b7F6g<K+=f]#f.45:^:Y=>CgOV:UZWaGb,E3c_@a
9f\6FR1e\&[N@fH;?e:@XARE.RM1=Q:2XECJAa3>e^f&dG,8-B,JNgX92HT=-gH[
Fg0.G/54HA#e::KS[8TXDH=G,FCRU[WJ&Z@LWF.[9&0+b:VfEJ/85^VN4EM]fRO^
Y)G&<2&g)H:NN;N&c5,M=)eM4R?C&R:[;Y1U3TM_#O8VS8b7__3S2A0?-E&.@1&1
UQ0\(=V,@>JfW0^\F2-A2T-H(69Dac)\)a2Z:W-/7H[\.+LB^>P]e&SH]Y/\E1SF
d^NUA&O;aT4+YV)AZ6M(OLE-(SCG.4^V?UWKMD.IX0F.]F.\_.R@ef<FNP^U/PHH
9JKJU-&,S:]:a^EPY77EYgSdB,9(B39BfR3b<(/Rb&WRM^#67D^S^JX[fE5gZ8_P
9S7PecCV:Z0T>dJ&EJ[P)Q&R\^V?Z;@T\UUWa58LgY6(5e&CI?@E=B/</g9#6+V[
5X_0HOROZ[aaPITMee+@+bcK2UMQf75J+a<=?Sc6SDQVgMFeYF@K1QLG^9LTEWRN
Q[FVL<)N^/P2N?R2+6^>OfR\8#f=P_S:4e3GC==W@ST8+O+DX;M2M+SV7?:JdOL&
VdG]b>TG&baNXCdG@+..POaPUZ5dDbQW.[X2b]/[A@bH4)/57]+9-&HZHW8Z=Y&Z
+F1?GBWb.#;W?,GGZ(S8e1c<3I?0T009>K)QV(Q,8+aK6L.(UBa+Mb-U]KTX-#WG
4f1ge:/Y+#/X:4DG?2b>5cJB/#fDM@0H#.JMVN1c;dS?cbHNZ>_f5Q=7,0;O1_Y9
W.-2Z:?F(?bH_5+g:DfZ+]&I7FUXCZWA-/(3I3+AH;Q?:A1#U31Kb6+51LYb7BUg
D490<.&d93,:3^bEB@Ya]D=PJ3@]f2Q1_KY-]7.-(Z=>@Ag4T<V+<47Fg#FSQ=gH
M]PV;BZSI7,0#.J3;V,W<[R/+J[7B=d<E:G(=::,PD,b\F6).-9)P3F+X<O<E<^:
A3+[>VTcgJ(-BQP]VZ63Qd1;D:VIeC(Ac.HC.[ZO+IR&ZBCPN9UI\a9^KQ?Ne@B]
C@O[07Y;\R#0-)6@^\QSdb)A4&^8GM.KR,5/7dTJ14dB8_#:,g6f&]@)c/6);L+N
def]VDC?#S1c[O,8P.O_,JBa0J3R&:,9B#=(EBHGZA;A55^+\6&c=RB3(M>)/eR\
N@e<]3@Y^-b0YVe:?^+S#KF7+VJ?g[G+:X.+/Z:\;P3:#-R(4@?(76O])I9ALC=_
6E]XHSc=Z,)31Mg,DE<W0?(D\IeTDV0P0gKIE8+1<JVRA>d??S+84f1S=Y[c7X-L
/XBA2^CGXI2;2g2_<KA^33EYWUV]41&&6@^-UL97A64JS\BT[Kb\,1a)4+f<LP0=
/PAHH,#)Gb#NBa49[=2ROgcg>W?FSJ/;gaD4Z[P.W#REdPZ-U)5PF-g[.?^PRG16
Wb7M_.E#DM0/500+[BJ(IKb<MNG)F#T,7^cZ,C3GH]>d>WG[=Pb:=PeT,aIJLe//
)15LCTX7OULQ9PY<C#(O36Wa?PKW^<Jf^XU[RVVAR\9#SDIF3.I/GE/=1PNN-U)G
4Ab85-O[VA9\E>CIFJ@C5L9+][S(ZT,VdU=<gK+D]CM_HaJ=P?<abHK@2TWYOF\J
UE21P>I1,&D:L0Tb-\O9+1F&<H0b&/(__RC=Y:&TEBZ&ZC(]L)0F,&48B.B+^DJX
=:.F40M[BX,U;dB15FVe.9[]gg[ZNZZE&5@(2eHYP[ad8V@^a@UQUX:]gGVTa),G
^<2/B)b6\G02&47P9I0^633a^XcfcOHJ/8?/H@N&#;:.UX4M)JZPdY&g-c+QfUX8
T_<;L5+fH3T2OfQc@.XW\^BAA&NNA0AI)/e)3;E,,6^M8_0;2ICF3TgT6@R4CcQZ
<T\&/F,1E9J>MMO7CBX?(2V7D?WJ1&5H&C;ALZ2A4/58&U<YB7F:^-,NU5F-6P-N
8&W8S/XC860dd)ITeU]M,bJ@KV7LTV..]@0N=11K5JK8[BJ/LGW_E;8Y_=FX08XE
Z&eH2L76,]Q4QHR6<DIdU72@.dFaI>G/N_#QNINW[?VGa2M@Ka7&Se.-J/1@\B\=
-0W60LI5J#OSR&-Ia+(J(EO)-M,9->^PEa+JAc0=C_?5B?<#a7(@?LGP-8RK;EY#
NYOd8(PYW)K84@Y.)Mc?E:SE?UHK.LRI6J4<)2MeTT\0aD&ERCAcTAW:WXFW>_W5
a.YA33gLZeNAT,;&Y)4-4P9a&V]]#>cd.K;QADS)N/NRG+)X64D<^:;@OUc=;7gC
.9T-R2C?^cb:3GfTUB-WM@6DNCbA3Wg@c@,]F#:1M/e__7(I[VZfP4@U[PUc4]6@
(^NbAJb7I:8VgeZ&3+)NQ&12fQ_N56O3,GQIHc@ND<?G^>T(-](G]B6EUKd;[?fM
1aUC0/M#67XR;J27bB+K_,D+/BfWELLN87WDSK1H2)Mf:a&NfO]E,/]Pa&:V-&M(
1,LYNJg4<#?a0S+.2^EgcU\L623,Qd;dBb1N&b>g0Uf<H)V9M0NZ=eZ.Y513JgT)
G?[CHdT^6GWWBX/e]QUMK1&9>54_fAVUfH45EF,NRag#0M9]_M=&V<3R\1#)Ff,6
7K;(&XLE.DVYIR_WQ..LP:b.?e[]AJU1,d.g(Gf42J\2Uf,>dbU0?;6CC:0._:&J
U?1#@[e0J+[4WVY2K&@T\#LK&T_WN^7)?I.b^4>68LPUQ+_bH_P1,GI2HFRf<X^Y
=\-;=F_c&O,G))_E0f/#gR=3;(CSZ)MO/IfEAK4V7EGaeXNc33PU2.5B:N8G8bO)
-6-4N&c21UW3C)c0#0LOP:S++,.)GTA[^JAR>]IGZ1[1NXfS/([,8F]V4ESbO/NC
)J+<K7L-)BVY)\L6_We#\3cac1[67dJO#\,8a)<g9=bcW:gJE=IAMa6J-5/XAS8E
5ddc4U3S7XTW)e2EVXAR9KVV5;L4)9U28^XQa-_QKEEJZ22+fPbIP>58/70<.,]1
4W>1F_G==-:17b_e[QGY?GU4d\-<a5Q8aO@_Ng:U58H\@cMI5VXZgU)TSWS4Z-#P
E<b;FgP9KFe06SU=E)D&J^&RI7D^d-AdgHV0NG4HDLP9Q3IQZ0WZ?Z)@#0Y7O6P4
FETLQ4+]aH-D.+5a4US,]ea-YG;g;VJTD.,R]KI9ObEZ1W4P&8&((CJKJ)FGF(GC
:5]F6fbPKaCc#ZJf8f?O2&<S<JD[X3f;2;gLQ8&QWcaLW@f8+)<-=T]OWSC-I_V0
^,EeR.(aS3XSMD@^VC_H)?aKd/#@J3>T@O-)(gK<CbQRfeI6RB4/P=AbgX#@g:UR
Z&[-_6D.If-^HdE4DU)a&;3Ib.F.Ya/O5]D5O.TQB@/<49fHQ9cSYZ>,/@D:N77C
2A^0KBBS7-U#]6.T#2cfcRCSaT?I0R9,/7^9H3I,G1JZ(X-MRM&^g[-D1[EGD9^<
Z<(KJ79MKNG&3fNVgFN\.WFA9EQYD2#BJR/6YK[AZ?[:F6]3KS_dQFfUb?[P><EU
BK<9b8=FQfIAQJ>LEI)CTBWeH.bH<3^I&5PPC@_e;NB5B^C5cY2Z)7aA8@2dQ>_c
?F3[3cA4F.,/DD^N/7c3We4=)Wf?T,T9H48S-9L#2)EX^NfgIP6aGK9B?KYEgBHZ
35O[/(8.GWSAFBA:5)#eC)#:f.edcUH(E0[^)C2e7FU?]5OZbR<ZEc>KRRR0T\eM
SfOg0f[OPN.DEe3#6ePO9.a[>b2da6g^[-M<f1KWeA/Q?TC,N9.?5S4-bB_dbe:[
@9\e[]S@Rac@QgKN,-67/gO_dd#5N18QAYe4J]4P<(9:Fb0AS_@_8G#c-<[2JE=,
I2\[E:DRJM;Y3LVGQ<Ka><(S[a?)&HP67#?PJPdIG@^F.2[WSSNYcZ(QSP#XY5RM
[dIS<V[eYZbX2Q;4\.2PdQ3ZO+:?5I?.<cPFI1#/[\5g7#aO\04YUUIYKK=W+7A^
ZEKe3AA,;Y&7K6;9.LKa];CKJ++e176>/9-cDXB/=4NMP=C(9ZI.;LObP(-cf3<X
PEHTb:0P>1C9HO>SV0aS^F>6.;Hf?/-7R5;8](?&e/<<c3&#6#:(R-@\J(4-I>9Q
g0Q_AC1P/\U4f2S-\2QYK61;URV\6&?d2+4K0JNaED8;:LPAW_EKV2T,T6EZZFO/
T\J6aKNXPDZ(],_NYET<)H(3X;(57@2](BT4F4@dGKKe(O)N#9L5TB9W2.J^LUQf
H4\:H<U9b@f7:FPecX+f;0TU?4>W?F[4<E&-2#^HIJ3_025?=[=O#ZYUKf&0Fa_F
G1baE)NdRb^GKOc&[K,,>Qe6&NYS6g?F?T.F+[SJ/)8#:F5MWAWAbH;H(Md:M]?c
8_QC4:;+<\G/VGY\ffC2\CX[+I6&J1gO@BUW.L<+B1aR9O\Y4Y&H5G:,g:W12OXA
0VTPN^7_07Z>3ag.<4CgBE_f_T;P>S@J?VE=R0B#&\1Ae4Q/D^7X_7@&SL<31;1V
BP7_?+:5Ce,&YfQZ]bGVd=/]J(&EE>9H(X3f_#Y0<CLc&K0_Y]Q@D4W2@8/6-cUb
T5-6)1ZUe(=R4A?GU[B&GA5^Ea>?4(bLEM\62SbJ.1V01aET@>L6CQ9bX6WdEY<;
8G@J&MKWf,IaO97.Gb-&.+@]?OOSR<6&6<E4]^A]^d0g,G)&449]5A,&-HQYZ9.=
T@eLgLEC\2[U6NdcJQ=Ke53IIRdFcG<fJPX2S-4^6b3V\,KMIdI#DR(ef:(X(c<7
XS>[F6C\:.K3I#=CcC1,]Y+:4=g=^P9+;IZ,.=Y&1;S^7-HG1@JYI,g@#3+D:+S/
HT&JT&@H#d_YT,#?L3(A2G6dbTXL?EP+:ef/^;?I7#]7[f@6)Y]&;8.30[fR3@)-
68&fAb2W,7Xg9,#1./cY2U#K-UZ=^X(ad5OCJJJ2Me<CI#V/-<5+641,_L#cEYYZ
OX<C+7@#+^7;0K2R1g\Bf9SU.0DCN2]4g>6ZP#CQd@G+c)+2>->C4+1-UbG/^-]_
HS)SLN#gONQ?7H.MP.ST&3C^2eEK+U^bd[-L<-9WFMRXN]1;^5bJ+=J,e[@=4,7g
Y(C1+6MO@)<_3:I.&LVQg^=DY60H[XR4W9[6]Wa/WeLX1JR,@Od^CU@+(ZN9RBF0
8=9NO3-<6ONgE&WZQ7^OA^?XOE4XI9(?\+<I;dMJ/Y^5V4PGRb^UEC2+A0P54GOe
6S.R;Ba0P>/YbWT&A6N)E2,PA<&M/M?fZU9,=f8[dTI9eM[=M.T>8#<&#b@CDKF2
H^W?L4:2=>.WT5R>K7e4Yf<WJf1,\Afd]5RB-5E/A&LQHLH^4MF<24B(eX=1[>c>
8db^b3O\5)>Cc^af\XF).?0ZgJMT)8/Sa0)UIRdWde16U](D+&gH+4g^&N[6O,R:
\L^,9Xa[PVggWBbD,gJZ5R=aTHDAR]80<??DT(d-(BNH,f7[2ZMc.L3eXNL)L;:K
GC-Y9<4AKM&G:5c<#@C8<B7c,dEZ)W86F#]ee]MBa.523+W39aBD&-@4Z(]_WG;>
5B7U((C,2DEH(GT^/WK(76_AL;c6gX1(46XC3^4fKIR)3R\7.Q&P-]JLANN/df+C
P/D0@,H=+4801?=NK2?#Va./KV&1Y8Y\&d^.T]>a<HX(1<T8E[H]Q82G&V8?5NQ0
S/Y+EE^C+dR=][(A?@UJg><JV95VDcR)Uf\S8QEe/2HBa^YBBa)[TfPK;W<,@c<D
:XCF/DQ@/.>T5Ca]Weca1G14_S3Tc]27db;BORJXRWRM)4DF#dNELHJ>\KN2FSW:
)FD:8FQC.G.+bBMYK+V]NaCDU_L=Wb+=(<?:dV]eVcD]/C+^JSAdQ>\FFGGc(9Pe
Ag1_=dTQ5deTbK+\RNOMUeHMY_Ed-LQdL4Ud3CKY=bJcH;I4J5,TOK0PU1)g9WEA
1FPHERg/^K1KeKgQ(R=d3--C?g4X[g_YHYb\A88XB?H<?6X4:Bg]3R93RQ\1VcR(
-Q5;WVa]=7Q5Zc<)<X-PM#V2,Zc@ED(2:gCX)2H-9fa#O#FG7FaP:6NE<)DKZ4=V
Q^6HK>(FCOI0T?+XI6=A#JUg>D@EUd)>?f=>SQNY=e3+_5.Agb:TfHI&37Oa_-;V
)]:QCT5>J:@4I)\H,X?LX:MOLbLeca5GNOY03=WG104:^UT)@P#aORJYDJN^N>bJ
b.]1(dO[1aM-NP8U.@dIRO3WG;?;JBa+N??XXIFS>3IV4K/KRK@)2ZSX0>I7>79C
T1C<FP+5Og4f_ENe.3aH[CP5N#S1UO<KBA1/IP1PEgSR==9V(FZNA&&1U05/,.?T
9/5]XL03N=BZaIWWR+H2@/e&?XHE:AMP5JG5JdN+fWL]dE39f>TP5CdM(V70Z>TQ
B(NB/Y[e=NFe5bX4e1P2\6L9OPc)XSU(=+?8XNbMRXUL1XG)#72ABT?eWA_&:]S(
)PJSYg/FNa(&Q/,GIVX;L4g<AXVXK382ES]3HaA97]:BLfEQ8WC;Y/f6E&/_ZRe,
JgZ;-T017KC(6&+GU0??05/)D;5D&fH6+S@DXTcODR#?69aN6_YN^P-1B8a#W[)S
Z?BG=bWIc(/)ZH&HY)-cDbU<U[6WQG/-bU:OHJIG.+&]O_ecVHa9K4.f_70)V+Z^
0<A_LY&#P++4N?-WWM>gGWUa@;YcWa531\ZO?Vfa_=#_J5TOBGX>4>^GQdBN#_cC
c:>+Ge3Bc<A]UdY7K\#B)RJDXEeP[,c/T7K2G2G2M3+aBU8M78A@\)e\^#FK^=ZP
M7Z\^+I]R55Y#GTGON_<fWU/DGeK4E>>5/dW]=e)IV4L86/<TTYIXR5+3MF6[?GM
=27YAdG+#^)L)eO]a<U?@(.BG=;JNb&^X[E@&3]c:.>aU-c3dY@d-B.O&4L&L;MW
3^[?+VOgSNJR/EaE[XTT>^)@@Z_)7L-Cge5Yab,:(FAg5=RTW.DV:YCI;)Z]K\4H
S/5\_G)Se<Q<f.N@1aaO48>WL5V>P1[DO\J^Y/M^NP_3?CWg3RO]Q[7Ef>bH>&86
O4^)3]\]Fa5]B<R1U?FDBQ]#AKFM,[NI?SBK+#A^eag:.N&FQBSLO::MHgI@Vc5/
0C8eg->2eI--(;7ZUMK9b4Y&9W5d>D5ER6=E_9]43)P=#)3Y(2_b:M[N_eQ]SZ0D
3K68GZW3AQU5XPAeP,?37L-cJ3P:J_+I19cDR_bLEAef@Ya>_afXKe.[[Z9[L0JD
MXa@,NdV-VIXIWU^8EUC.&&Ie&^2E:.eXOfaBJf5]P]9+QA(4TgNBZ9+L3/IWFTN
Q94Bb/Kb9)_8A._MQdc)8RSLC.N/4X2H(>A]eC^/,XAV5ODVIX/[KOCS@VKTE9+?
SS3DH49NNU4<G\+IOZO0X)<6-98LK?bc/IbJ3&@?W:0Dd9S+@=E.838[0OcU9EP5
0X?O#8Y_b39/VdeZ+-HO_eL,W4O671>:&>1OM6cbcW:586F09AW\0C+5=;1SS/OF
^Ag2B#DST)f:2c)BfU^(45.[DcK4D8?GUOU^(=B)N,cU6)]BeXG@cY[,SbGICXe@
)8^[4:X/7\=,0I61YE/2H[DLN/+MHc71?fQQ=HX^WJLAI[HO84Egg=^;6SSg8U&W
7QKH_O&1KcaJ;@VZ>#a36>\;gTAfF.3O]QUQc<RGF,L#L1=34U\73\XPX2Eg@B#1
:dZ(fRSPgPb)&,G#D]b1-OSHa+3g<#(U^e2L1M\6F16V:D]H1,\bNV+:8FAZb[6Q
e-/Z<QT5;M1K<:AT1cF]ZGa7(c[?WH-/2Ha#H2aLMQfef>J9YOSa-K:W5;A7B5d-
cEJ^KT[-+d@f5b?2WB007.BL-D=GEI@U5]FMV(=J:96b]Z@GGL5^/<cT6@1g@]YX
d3_NPZBfB]P4f3=Re7GP2&RH9//F2V/J&V0SDg.:/dC^9IPXQdK)AWPRc/+N>\Mb
OUc+B(9;GPSBFST;AeA(H@c&:R3YaTdPd\O4QUF<8P()+G)-&dCE@[^gK[AFXZ+E
UQQf5E4T3L<B^O/EUSHV@bFTKfcK;#-.9Wg>d@IH&3_@(C0NW]J(-Z&81?Q^91IP
[eP)bdAF+8Q6P,Nd,_O(Y\-3fP48b;V4]c\O]@M:VMR1-MP=8aT@:;TIYbPZ-BcL
V2>XZ9N=G]_2SPVeW\6D@OQE.J,dFI(G&-4LDFJZ93[E(eg3,<MI@L)P&#Y,_3/R
/B@)>W\(,;2JK7Y9cd3[4gHLZ5<<9.>#@R+5WdTFLZUdHG(g1V1@H(JSAU2Z[O8e
S)d75Afe4dZ3^ZHJP75_f<[M:D5@,fD8)U<7SL/8>56(3Nd05R14NPG9JKONA@6@
CYV&MI/Ud4,I-DggW,b@/O+R&]O,VY\B_a13=D:_-ZBOL.MU=RAS(e/Lc@FP,FQC
c;8GG#1R@@5N8^E^c+19c5]IOM9GcUJNB)Q-c0&>^ILG_61Xc/ac=bd=b6XgeV[X
QX^>G@f7A(bDF\(HCG,_.YS7bVJ[SaQ[Y96<+NaM])1G<UDW^1,fGNL3Ua]HNW2<
4H1ae0.6E4Ug9Q#ODggdX).Z>3fS)dNP()#39E_W4U]43/MQMD1(5943N2cY+0?-
?f]:g-bb?##dacbeUb^:C]6Y7D[FfTaSUb7OE3)e\#O,1?bQ)&(BLI-.;=56>ZO+
1=9baL^Z>-NJ=MEY<3:_UI5?^CHdg0OTHQDda_F);A=<P[GN\d02N&5FK_GH^;AE
HdfFBDO7=>:ZAcQgJ2.QMPO-gU7)I.9b59JC3\QMR5aW-/UEY+,a-JBFgMOG]-Q/
R:S1Y.7/0GHX]J+N42^&CN8Vf\2RMR5bX[FE<8H]:9PLNZ3I-[872b)eOGO,Bc[5
^RQUOcGdZ<)>NB;,@:2^QY,_OFL,UZW5698\XI;?E;&<I7[Y&33Y7A_:^?3[Qc@P
+e35[^YF<6J(I<dT?BV4^<]fE\Y@IcI(0BDNZa]e]ffIX:G<FORHJ4P<:ZHV7ffT
A3\IKE&&WP_<K++eG,97A[5KbG4&^)6(Q3)>fc6)9CDXFgRU+-3^>N^5Y;,J<AgS
8T4_ZJCB,8-BXUSXA>VK<f6Y]_5K5#G,UU0QgD#T]&cfZ(2Xe-D.YNa<dgD#8496
>b^7F)(V.9dQ@>afXSG\5eS&U]1;?D3T])^NMbY;7;19MMLQQf[EYbdV9&60OMJ+
F&.E2NA5Da)MYESZ?4M#YC3EaMe@B0EL6I53VQ<B_eE6WJ@1F0P^;V71Ba-+f<VI
.U#Z);/6SDUFY+W9]b(EaGY6:V)FO-CKCM;W/WOP9a^6>,,>;?]6e#a>Ua7Pac[[
:0)-T]DfUO[c<2T@-DYQf;KH8@O(?#=b&\f=4DFgXYEETYW=daX^(c)M+E+K8cYQ
&ebgOH8G\)WK4X?gf0F+T&CU_T#d[O<FQd438S:?VT@K(R9O#].M[A3WA^SB-??H
A1?4-,NYO_2NfDX8OdIJ^c+J[&,3V>.e5:R?EP;[f\T)=cV[?B45?d4<6QGJA?P8
.2LgQYU12+)N6e_6)R1>g:bV71LWcMd0Q\92[9A9]C68).TDSLZ@L?+O@WZe-;.X
KXR/3^<89JT=J<EK8\>+Sd06?dTV]QdZZB+#,C70O/DEU)#Z9cf^++[&15U][(N1
bgY]C?9P)B70RGZ=6/33CKN@dcgH(^[T?Ta1PecG-0TU2L37ff(IBR?DG\R,><.G
TJ(N_XVIEZLNS[Q9e^]PI70ea,R\&H2^&)WHTfZBc3(S7@J0+JHd.,6VUE#SF)&d
6HHaZZX5H1:.80ad)>R4JM5FB_A:C]H+E/,FG3eBN80Xc]FBA9f_Oe4_7\=78GD+
H:1348FaF/>-fW:)=<0fc>d/7Xge_X=L^QIW0#=#M61DY29]15KbDBV16+0(N5Ac
7]>g:9Z:,X8F4F-GgA-Q:[VX(T2K=2IF_fa]2dTKLVR-fC&XW)V6CXTa9>31X+14
,FHPE3E^C[T.KCS8EG[8Y>[IC:3.>e0?;NbV;L9gaQ63>[#9_1K598c7JFHXCBcW
0ZX.UWNcdP#e;(MEED0UO)RN\+2.;TBI-0X?#[#1FOb934ZXFE-bAX]BTE8MMH?/
:E5&QX4Q/aT#GPQ8;,cT=^:V?[\P>6YCAE9,BMNG,:8V.U8<fcdA5g=gSP8LOZ<M
>3Q\1+XB0Pe4/KeTL8=Nd(-LaZN648LF7LO^[O#Y#Ee+(?K/b8Rd.Q8^HJHG/@GF
NV.Tg3>HTX]58Z=ZXISM.AHA.7GB-HN1GZ,ggFC:9R>X]7I,O^,,U<:;,7PY8D<)
U6Kd,e_>[,\T>FWaINVA;ZQLTL[92X.GJNGQ:AZcA(2C)[;g7Wf/ZfSSC2QXOR0P
7C<P>aZ<&WG7PPgZ#?.:RKJCCFZ;AgZe,S>4JE:@Qg522@-H9<KfYK=GfY_SJ,)g
1c/YD(QFK+FgC4f&HZ6UI34LRQ>L5]]+(-\a3?eE;1VP-/:_GGRg00g/Y+SY8TSZ
K78OIZaE@52<)GJ7?T7W]1XV5&W>X#Ed^C;@:8AHcV)0Wf:())(\YG8+ZWaG5?.L
\KK023KD=>b@V/&4c2[S8RDgaI93CB9S;)RX#YQH3Ff/Q)L17TDOQ]b._a:I+Id-
A9&3Y;4AE\X:)I4;A62@UC#KVKAK\JB>N5XTL@3gDW=-M7-e-<Z24=I93[@b#<0\
>A6)<3&:]7-#@WMR?C6;)2S8gY.=<OJ>MU+.Pg0M+#^L;N/ea7R8GYZ1_>BL_UWF
637E4LFENMN/ebI(8^<#_]BVJ_1c#cEW=4_O^g.MQNfXX85Y;OaOJ8HZ;_GPF(RN
f];FdNSK_YWf6U.Ee1+4:@<\<(+L1?8,=+RMdI7@2U_.gBd\cFZDg.9B=5:gXB.7
Nd:,dB[P/cN+O(R/M64UV1<0=.g:.WV#KX4R.Z1[WXSNI32443E.a036/+b/BY97
XQMed<.8?L3FaV-MTT^(BTVOOLRZG^2MGP&^>:0/FB>R,9#?JNMB,J[(+K12VPC1
#8:0X\GYLa_RBRFHNR<N;Nd:g;+INF4;N\);dWA59[PZSM57gH6X:2G^WCd^/7gO
b[=F-E04&)@@b9R@LBg>NUO#fUaJ\2&)fA6f0NE6XC0W\0;bTE0._H7V)S/[2edH
cD:ZUA_[Oa1<R,CS3>g(D1O3IE#1&5,0;9705)^?9GbcTf/PeeR^6-I4AZ^&6_?4
POYMJ40H_Q[5)C2<N>XZ^bWDYRf9<&?CQ?[R2a30=cYO6V+VFf#;II;DH5(0E:P^
<65.+RMF_IY^cMQa#Z9;eYT9=6CW.[K]68@_7POX,9]f?L;^c@5dXd-X\;UQE^Hg
NQ8G0FWf<S^X,U6^7Jg(VXNUeSP+EB^9fO])Le;2QZ?PC[AD@e-(/6:JgG<F5d]R
;ZX^6HZaTDcbWY_)1;A@G?TX+-CH<&97+M@3Pe^UbWZ+#a_b&_/OF4R#)AYgHF3_
=8ZN.:[,M\)L6LNd@dU(I#@;[1-H,X8a\>Y/XV9B)(AJ)7NPaW)AJREMRg<Cc[H>
]4+f2BfCf^<=GBVXW&gQ&8#XT)JAJQE-_JP@&\b^eL^MQ^3FU&aQR@ZF&5__JL];
b8NJa16=b5N7=Z=bGa_0\AO3\PU/+?b_8fJ3[89?eSOQc.)1JJWS2MaNJZ4GU\K,
Ga6Gbb^e)376,LSd&\,R8U):7O=O?6YF0g=JNO]3#W->;M?AMcU[K<D/9QA3FF49
116OJ^5R3.?9Z7TfOX^DV\g6Ce#L#]GHR)^f_;fE2Je&4H613AR<I6[CeI+e>+8X
<]EZ>dPaAF2?7@/E(R5BH(c8b&E?Q-^CA:fXe@beRV1&,F3?)#=T@SfT\?f2\7>b
e^N0^-;I&[<;UQUTZ&0c\G;;XNTKcC6FR)F\Q1\Cb50CAb#[.U7[]?/)C\T&(67G
1fECLAYQVX(,YC4OEX@]-]cdD(X\+af.#\49.</7a?D][H(0D7cQTbM[8PUFeKFD
1K^+ddB]We&IHgfR\])]aLEKPBA4^=ORI84+FNIJ#OLR6B6>8TE#De:+K7UU>^GI
949_.SRK:d&XQ?W0NQ29W]]YII;)]P7@M32QYMAA[-GO)Z[5(LO)+YBV,QG.WM:F
-A6(4W;gVXXD5?7L]c>)SVb#WgAM/T/dM44XXHgg.<7;B73]L/cO(K2OCDe[TR+B
bE,cYgX+@,TTG#KSQfK==Z,4=@IcYV&8V&Z99#9K499/]W^11X><3;G3.eM/+J>G
6:/<-^XfTPe1W1WM)Y12gWFB(AI.TGf06FfF^+R9(#gaaQeZ(DXBQ[,gB;L@W0VR
RZ91JD_6=597W#)8#4(?BNU5?QM[A_5:GW_dK1a&:-@GNDf(QC(<JD^9ZGGX^3S\
:gNH4/2TS;TRO7^geCCM0662a4f5.XHGK#De<-\96O9SVe4>(>[2[TR:LCcO[Y)=
bTJ53VNE8fF]4D_G\R,5f@X=Hb+Y^F7;835D/0CJ)M2M]O0;0Eb9</@Tc]64^<K0
G0F=egb(K6M2TE=gZcF-]2g2R2HWFP7OGZU80[Z[)E1N19cKLcVEDZeIA4X;IX#8
@2BA=g5:>Qa@#;FV>eRP;SH1cb)IeNXI@:@DP]TI#U37L2?ZQaS?#V]R0\OK59HU
7,OVKX:aP:PaT9R]77^AXB>U3/..:ILNZY_;J9F>0dE@IURPJH_)SQAMV:.c#X\C
A?YU_@BD2d-;\F2fP.J1AI9ZT>[Z3&ZJG9<4EdR8fH<J@Z9H&7Je\[?g?BRFW=<_
=FA.6^5aVW(?:&>W<2Z.36RMIKffF75J.eg=6]B0WdTDP5RQQX1+aYY8(3AZcNa9
d)B=?dP7);Bgg&AIN;+OTaEB9#6Z[)0_=Y)XM1&^&=E_H#_GeBQCB:XHK,?9Wc;f
MSa8:He6^D^O@]Ob0.a0C(3+)?YdXT.9We[\]dYF,/bF\477d[AVC:PN>4ZU=)9R
[/?L=+?f3KKT>2;PWb&a0aagF/MPe#K?G?V;J4TSH<8D&(3S1d09\[)b:L78B0G)
)Z?E,.-/LH2WD/e1&3BZ)f&3R;USO667G)Mee.ON#P+O04?XGNd1Zad\H-AUJ(GU
W+,501aaSFGK>fN4b@@e&11W?R^6fZ4(=\MNSF>C]e.K/dcW335/,+VY5G0AEZL(
=a4dY-_cB=f4ZT1_)(Ve4BZ8P36]#&]\aO3X5SX)33a4R;)_;IFCV[/5=6Q5N-Rc
RHVZ(]Be;S^)LH9/>=H?[;L4JdYI+)7^:[a3[fO;6g-Vdb:[,Wbg=O3dLecKH12N
&g2?WAQ\Z-,O-YONK7NSD8#AJOe5MYMVO?0g>-,IfGGC?]e]#8VOG,KADPMWGY.Z
<G\WI[-]YZPTYf1&1V@FXCR>DN&N6HVYLJP,Q]_L3/f:^XP,&^b0Q,6ec&6[WOP#
eDI#BN+??Tb?G3^/2G;Tg6d3S2d6CH\]d(/B[CGe+c1G<]b-R@2gH0E6ZK<WRY,e
+B[EJBE=.[Md-59GJ.:,=2#[@17NQ[HFI>6VC;V)-g3,CN3+B/QCM+?89VBQO:K\
1dEL#K^.JA]Y#50adM)e=:@bHNZ5;OdTBBN>=7]6G]5:Z1\9PGZTQL,[(O5V;V12
77CBUe<>fG_7P@cD\U0&MOVB\&FH&L=_>Q)gWP7YY9:,TDHOA(,3J)YPV#\<H8_0
C@5R.2?TcYe\ZK5^UXOB=^EZ)4/DCGd;MFLH_JY3K&VR&N?1G<MSPUY1I5E\-Z2.
W7_I^1M+O<S4eM3UeY0#f?]J#Aa:\3_23fUI]O3(IS.NG;gHX:LRX8DKCI5/BAKZ
V>O[-W+#4R#3.>dI0Y9SSG&I6ZF:K7UCX6ZIZP3747a[b9,QNH+;g5)M,,/.9abW
/W[+a77R1@T\P<8Ae^GSKf);d08Zg/DcM61DMK9Xdd+IO#]<?M27V/TWQbe;cM\\
N+5;4:MOQ.SQIFa4#,;:R_2T6&a[cb\WOTM3YR]GR-H3WBNBebK._e_CL8\1E.K6
_4UPY2]II_/LL:Y2A]V2Z@X([<OQ:238#Ld@T[]fF&R-URfgE<d,V4B7]YWd#FTN
D/f@+DYGJALa2dZPJ?2_gA:d6YRIPQHa+F<(->7BZ2FF\/4cP\79(BFRY5]HLgc4
X=KE(E22UE(#.^-1>Ja(AfUd8J+2^?J&:.\g7=9#JOSL\,MXXEPcc<YJ<fXe\@L/
3V.\=RW,]TE>]2O?.H+5DacVg)#M26\EMffSfR3J0Rd.\&M@CO>@2E^bd5.d.@H@
B8X&\cH90e/U9]_VOZ_=76>]ZM9-0]e.F+C1/UASfD(RC=bS+WR<48bSR.)eb^P^
fd0T@,(=6P.WV3W1:(&59^Q,e4T5_7AD]S3BMWN?F,N-WSJS,@DeMf.d4OfFJ:VQ
>7QE_A)F[7-1EY]UbD8MR9.J-CS,T2B]\+>?B-2Ye8+\8-A0e)D&KSd\O)+2PNL.
b:>V=Ugfa_/6Y[;UDg;.-O4&K^RN<)I]-6LVZ?V&QP996/#^TI[8A50U(UQb#fK6
P3OR+Z1MIWXAT9+dc8g5/JR_9U\PU(O..IcJ-3)H,8^E(:8U-89#EP._5<gfNBNF
O,NWdadHUAG_.Z^eK9H>A/-PN9Hf/)3Z.:,C@Z5#&fT)>L-2;0\/U03>NO/EdI.&
F.UQEe#YQOY8CWXVO6CeYYcJE,Q-E.N1g#Y57HN:a;e=eP5RXGPg(V;IX5#)]<HK
CP4.VM\ZH)S9EBGXf;;D65M861BBcDcR4g,E32fdRXb;CCA#AU,@aDKZ3/XR+XP#
f1)-_+gLMX7fg-M_XWd71OL\P7QNR0V;9c9aZH9R-a9C<=TZU.^_be3530<dFI\(
2-JCMc^7a<OHV+CJ_I5M]56,cLAcD)3TW&e=NQI\RI]MMRM_(3KQHf.JS1>Z\L&?
L2,,=f,e,M;7CI4=[(b0TWZ>Y#T(OO3ZgW;>FHf)bQ[XM&=UJAOe:99.U;9ZH]5_
X,f7BKc5C,d+\:APcK,e,ICaUSQ(E63?AL(+M:fDg4,-e#7F5,ZDEMa78I1V[BU(
G[Y:ZHg7>W.E1aWeXN4#\AXV@D.(.#]WR5g]Mb0S3J^g>45TVXgQ^I_MLgXFO_:(
Y@)b]=e;Ze&aAMgGK-E?EOI1cca5a.7INfJSDf2Y-3>PJM3_Y>A75MD]^gXe?K3W
^DR-[]H8<:D;@UK7N^eTP/b)0BD3d?4PN8^?#Q+.c<ga5a+CGJ(N[MI2NNI,G[HC
7][O58IY]2gV[(9V-Pf>b,FUAAM.CM,c#>1K0.4K4P8@Vgc9deR.(Z1(B)bND@:N
#]5cBcC^)K_.Z7X;AZT=N89L-:_U;?1=MM>=DIb+^6L_b^K9RL@D\Gg[QSbL6fb_
#,A@9]cR(4SM\@5&4CB0g;[]g43T4<;MH1+>5:<+LRQ]4L95^4:7,(_#Y)&(9X--
G6L_Y6Y04,N<4:@?-?N<N>(GfaG?G+.02AVC6Fcd?W4a5IN(B3cS/Ob7[Z,Fa4[d
[OEH2:0<g9/,U?GP9GdK?gENK_MV@VP>(XZTbQ,gOSJN+/T_g3[gLWOM]CD5KXVf
>Z;JfY)<dS0/[WL)=<5.SX=,Qc(DLQ[H4)QaVLd3dSdcAAQTKa]UDc]+4_]bQFgZ
WB(0\PQ<B=.1<XH/MO/YS-#>OSS)^??d=&XD#WO@3S8f:d4R5Se5I:B-@3P[<#Xf
c)=?LJ(KfVDd38)-a\(J?,dR]-SU::c4DB8EX7b=8)/O0H6_3-K6LY+XG#g9B[[@
N;)OU^Y+&<J;d1UJMRDB<Zb@>I<>(6KfQ5d&Q\Ze)gEXeP_Y=.A>,IXD\>&:b]J<
+,D<T0,+4@C:Y0f^R;.-cd+QRO9KP]?+PJ?B0JL[bIf@:L]=M<cA/\2g>cc8cfc_
32<PB\C4+65E9Ted&XVMWZUONLYUR1W4IBK68(FN@SO5>+dLe^C^LQPPL>]bGgGW
3S3>.\;4)6XYW::LI;5SOYa0da/<-F#:B^Q8G5B;H-SEU<Oc_CWb29U=1>Q[_48)
Ae>X^;IB=@0c<202gHC=DgcdOd^YJL=K84;\WKC060SH9L<1A/:SB\_T29663TS/
Jfe^)(CZN8NDGOg16TU_^>65-8C66<QcTPd(;6L/O/>/g5=;gfKB[T<:>\7V(Nd-
9>&S+a38@414ZafH,d,EX-VU8U5:IEQZ,aB4SeZP/;3Vg2PH((I2X?;[/#aU)&Z]
5^Na)bY6Nef&6?</W8-Z+>J)Q4YD=g+LPdIS[C5\#^+32RMIY[@BIDH]S9b+0D^?
/>JVD;2#ddTJK4PYH+,MP]_P08bgdLSBOS4P]Y#/L?U4/e3MgOCaUASgO9gZ>5A0
C]WO1g.56dK9P5?Yg;976R_THQ,8R:Wg&3JU.,.DE(E:V+=N\-1D\][.T/,c_RAM
_;P)]7](AWFRCQ,]>7L?+cVH?+-OeKLX;V[RTJE;@dQ7HZT+gag3S?A+3_49LW4\
?JHG[:<W#UXD3-_=Uff.,OOHWDZd/MMgMMP[JJ#6X;5ReQL\8cB.14>XDHVX2dQ#
dEIC/ee[OK[,2,bE630]YJaT3\L2cKS_S<5WJ4A)OfYZ4;CZTL4bGPd4TYe)<UU3
0E#91[d-A84fUK-I7PBD>?c6(QUBaG+NJ:?\Cd@K@Q=KXVVEfB+=F+_9cFQMD-_Y
O7bSf7>Jbg<R[DDW@AgIUFgd=:BIRE&11R=RBR-&OM3Uf1F?FV5@FOF0XQT&E6g?
1_2,G0S:GXFeX?WB86CZXB/<;ZW)Y[:KHD7LAOWH(,@_X37OZ&S8-I?4M@XZZ1Sg
[[6_,JX99[N(c+dbY-V-XJ@^X)?]A+gPI?aS/K(2GZEf-;ZNO25?KS__U1C;B5R>
7M(P(ScYT>E1/6C2#KF\L6]/0\g987OHU[DTNUT5c<E/VYU+EEAH=KCB6LCfTX,T
@gOe/f]<)&13eZ;<QXd]MQ0SC+D\^3Yb#0fd0GFO,)B\2YbZ)3SLAB1N0LNTGc1S
=-<./AEOX4UV[KOEP;OQB388GQ7dHGdccW::7L65V;3,_J@IOGMGA8aY4>@ZdgI^
:;Md\fdU\f.XQ2Z+RFN5-,c)LBOOB[30NINJ_c:VQ8[T);D>+6b953Q+-,_E_)Kc
18Kd7LW\L\acR9:<DHWbNAb-&(5H,d#CRRba&8<>1X=1E(O=,B2E4SVP:E5YP6/<
a&):)4)VQ:Y:OM752[eMP2eF^Fc\+8-RX:YGg@56L)7NE>J6CM^5?V62Y2#U1_PP
eQ<Dg(-D2OI4;7SQX2BdPD3fTDA07SEbg)daa,Z.9GVS7g)A2@4L?W;;SXV.L=^&
JbM-I@NFb4F8(dI,267UU(TAS;2[E1>(F-#B4PV6]9&M[>-Y60^O<VdVTU+X=Y9_
dS<@P4_I.c0Na_\F7_)56\9)&0a#]bN\BgfcCWEKbX-U(<FGKOFMW,CPT4ZH]2O<
E#eb#ObE>,e^D1OJaQf_+[A3F&>,4f4.CI0/QGKX5=ba:IP2NXR<I\>0HOEOg9Rb
-9VN-K9Z?UM\PI8VUeRH]T(B2Ffda]VYY2WP_P4?76>RfE:U6=OddU;&]Z.&3TA?
MG;55L0/S:5\Y8/H8B&,Z[<#A2Q\QKEUZg/VW<&2<4F7ge.ESDA?V@;X_/\a^?<d
4X57U;^AOX4<K_-QPYMGV35\+FD&bJR)<RKPMgOf8Cg=A_A/HZ-)Pe?Q[?b2:=B?
=;[@AaFaV=N4Ofg:#AeIdJ<d5c3b0MET^MAQ?G/B1+VA9?^a;ERg#IdP3a7Xc3Z0
6fb<4g7QQ&EIEE,a]S,V^]WC9S_.,YQC7-+[ff@-FK&]eUB_B=74U7aA.?3gQ.J@
SXLO,:LUI/8_8aLU&HN0SS_EE7NG^b^e4JaYJ7f?S>]fa17-PMa>TF]-:Ia\OG5O
\QX&AINKVWO=+LY;>HZc1W3g\E1CMVTg674MEOR=B>1][fPF,J5VcF<52(I<XWeO
ZPXH6A54_90A(\BM6TC8L=VIKT1f6VDD((K@=dC)K;V2BRK#dFQdS.#(&MK]5^D]
Q:\[d[?2Ee0L\Mc[K2eA=3^:/+K#H/-<4TE>ZcD<HcNbaQQfL#UTaA9<Yf[H)=;M
Sf7J1X/S@dO-WS<IbEUe&AVO?ZOKP1?:Q)<^g;E1?M^^3THDa]Z)4^:f6G0/848c
MPHSYZ+W1_[^HWMT)-_B&D<>6I<B-+?7IDU2^a4#d^RJU/f]QA+I]Kb++bS;CbLB
BN8.7L4ebE@FPRUWDR_GYbM_CMFYe5>+9/X=?X2C^(#QV^9Q)?4L&=].\68,-HV2
Y\O()UU;ecCRbF.gac\J:)?=D7F\P\O9-7A+XP7>[[3>G5H35-e7-Gf&55@d+bb<
b)+X)+MY:Ig/T>bB9(4bAb#8S9Vb,+cK6:Xe-f1NZ,RBM+b>)Q6cAgJ5Z3X.EEf/
2AGLE8/(X>#db6cTC[K.)ZDaU4cUaP8J;4#d>+f6I>(O0c[_cOF[^_7KGdSD>:.&
4=DOHcWb<=;L?6+[I0#=?KZ9]DF7c>6?BA(JOA7c2@He&RWV.T<F:B\ZU(&Q/;\D
3^)d]?U+/T0LAZc4SCZbYPZPEW0^7C63/a#U5N(bI<24Q5IB[HQd+)ULAgT5:@;O
A6SHI>U/:dY>91[47@+AJ]-:RBJ:+5M]2\AF)GP,62/;1c0]<]QV+XTf-_J&[N0c
:cd;/:c99b8X#OVHd3K024MD)A_e??HJAS3(/+<G,#BXWR[UEX6W4+/]G>ebX3Lb
Z493RS9b;#E:PdUB.:0T<FYOFY&:\#)/0QMZ-EM,e5f/R3]<],Ab-KHXJ08K&+E:
7NdMJ-0Maa,gTF5/,<1YUSA[::3QD(]D5M6dT;7SE5#:4=?8Y?K04\U^:8B)?0-;
b1SK^@\LV/&^X2=ZT=e0E_GA,R9^/afD8YZ6J2]_KHMX:Z)W;aJ_XF]V\QJa:@NT
,Q8aED_J\HYAPC7H)Z:JC5,+,,1O/2?W_,M)7P:3)C#8<gRXbYH&Yg08.Y;IZ4P@
FRI)SFTXH90T4e\,UbZ=<QdG<e9+-8T@bG@8=3C9R?e<f3AfW=:J:FXY+J;K&)_^
0HISDC72PD6&__22KG:WFZ#JM]Ig/_6d+DY6CcB@L3E@+XVM/YFZ:KG(.\_#\L3?
FLc]QbgLUb<1aY7USFHMGGQWd(_]3,0eQc=T)_7KV0,OEOW;:/\BVe0GdJYdVfE]
Y0@d.&6>c\G@B:;\>0B&3AL,c8#I8TI)@(9L:K3+g^G2[;f\_)_6C#IGF_5VUT?L
UFEMY6D\=+KAL7)b7[W+\@PPc&-OR\DG^.3APDb>:Y_-CCg-R@<fc^g(RABJMW1K
N,cYG94[5#V,O?1/Q-E72^:Ua0D4U_:0/ML23DP//a+ae#7_QP]<@9f2PBQZ4X:Z
Q3Bcaf[8-\1G6<>]-bB[,D#Z+cO](BL/:6cZ=#JLe\RPf\T?.=;fV75^GP>^fcKC
(Z.)8X3)ZaSMCA_F)(@3?Rba&[R5/fcb-:<RO4949Z\>bT/<b@_Wd>)cS]C^C&J:
Q1M9_cZGMDTgVRHIa]aUDLbVEKC_@L-[Y<PMde+H27^D#A&agBVC2TYZ@&VS++=3
H/VI&gC7gZQE(+^FOZ.X^@<1^eZ02S:/R\,F\g4dFg1P0\<H9W-VaRA^c80#-O59
N08_;FIHG?1W<.V6KdK[)gIQ=NAG=1_ZI/\aAebf4YL@+W?6Jg,9W<9\J,<NJL_-
9R5aH^\4<^IaL-+05b22d^ZS:<V^OIe@?V67W#J_\11,1.BP1/H<G@Y-[.;YG._A
BTUQN1e?E&@)P8d5)3ZVf,D1?>ZWgN1g;QOFF(N/V#R\\1BYf:3X1N-AeHX(M&Eb
K0BNP9Y[^@8gUG(N]YK2DUS++2R</;PVCU2N&QYR[5,EfI1UO<]U@WA<+LE:TX3D
X4c^]eO_TV=I&>WNL)gD90S6<#/O(b5JU/&DF3[=9C^O]X,K1SV6;eSU<GH[>#@?
0[>c@@^LM-#+P?)OTJI-EP;C7/PgbK]d<@21IW8gQ\L-^8F^MdV8=_75=cAW;7H)
6V89E)PfCZPg7A__c.bVEQ.ZF8e^3]VGQSPe6V91V]O&O;O73FT6O/+<AN6E?BE9
UK8dD.MG5NQg12>.>6[f.S07b,6;V:SA2=,McHX4)HG2+HGe>c\G9aggZ>/D4+,_
65d8Kc]-=5T1;b?:[K[D57a(E346IJWD#(],,4ef:X^VPIQKU0MURgfE+]b(DM]N
Q&_G@F18:KLb_9S;FV+KN&-YL@Y3&-8Q1N<,ONM._dG,_6<XICSCA=I^D<:XBfbQ
2?S<f=L)VWXE?00D9C<,V?HaO3+I(0,f(,D?WG^:E@6cg;+X.TI,a.;F\09Pd8@O
L+;XG5EGTSPbbZ-cGO8H8Rbb[VVU,T^JKG@T8]#22[;,W;04,GDE69_J35acAP-_
TP4YM2da0Z0/dYP_WEDSK1#:QY:UYLKSNUN.WNVXGd<7>#dCNe-.4bgDHC4<MK.,
0Y62\:(+WRHZ_;.JBB;>\RU2TQD#e912Y7EXHVZ(0BT@I/Rb(+VV-E\C11;#\UQN
\7T@.66_F>PaH@\3Q/>GgNFW3=X^EC\e,]#ZNQ?78E3\<[SZC0/deJTO-\Ic2+6,
0U,E_98V5Z>\f2ZVZ=OW-Ldc22=<XDHE+[\]O..RdIDSMLQDXOXQ9^1?;HW8WI<0
L.(Z]+6F@DX&c?@e66.Wb8/4_73J<?<;&TJA1U9QJ?TbdCbRMU212gdS>N/C2I(T
.9g0_]F93PNfIaDe\M(Xe6O@Lf=X/O72)-4B/S>:;M3W5VZ/0#0@HGWZ(TLTC]\c
/KPB0+^5W7A5]>cW96Cg=DY@HeM[3\4E-H616[E.UKQF(F>S77G<X>[3L8>OCFe+
9+DI0D^X^NDQ9C)\d3[,BU39FO(Qd=&-Z_43-OV,:53EG]G33U08Z398HbR)Q>V0
e^_?L?QLZVYCOWZ<>>d3:GI0-L_ELMUJ[=GEKD<4WIX7Lc[#7]JJ8ZUPe<20L,HV
/>4[dXaaT]-e5<CADLZ=Tf[GfU(N<CU<c?-@#Ag&V[W/A/aaZQ:O0SbBIc08LFZ\
M:,@@bDYEC?.?95-IS-d7:b\:A7,0DN^DCTdKV;NRV6Yb3MF;JG@g0C9+5VDC[ae
d1TVB:@^.D/XRV6+QWb7,J=IZZHbEZT_//c>;:J9ND\WU@#?[KQ&_#H)PfL+>bJ/
VfF]D>K4[D4fPdZS>2c4^EXe>O./[QdgYdCDB?,C]XA6MF]])4^5bLDI+UVaG>Kc
aHDUE(3;1X1LgL;Ed5;55>G];XceQ;,>:1D&_F\#+6KZe5AU?g4<G7LRKfGWES,+
M-\<&LB[G.T,IYZC+I@EE(XTd+U\>^B/[BE?_Z>T;1bX1e=f-5,?3CEN+2<RC8#U
.0K.Z,]7Z0gR;UG]66@M]53;,^2;5\J)4W]@e8L8Z+5F#BegZ8KNK(#+R^-\YP)C
[71f#9(+fB-BC<dVKcMRZ;B>>N>]f3CF+XFIFSH<--UJJ(g8H_)Zd)e(2fB5Q>57
LBgLDOV@7SRTP1+V<-<=/fYf8M[SYYQB.87IbRAH/F?4.0<F,<JJPc0-F8FFgH-S
#8>R_]);Rb6YZ7GO6&#2dEAgG1JT(ffgT8,9L\+;S;eA2Q201)@W]3c._<0ZU55]
DO=Y)eaT<N]>DKf;L;?Z&28LXecY&D)D8-_JAe&KQV.Q_D)a=aS./2Zg0DW&T]-[
fW7CM?I+NM5;POPW-N1I+Q8<T0OVb-B@9@1\UK(F-6_YSP49D,OD-;8_29UDG1X)
\@bL#Qc0>>FC>>KD+0))-T6Y+a)V01FR73;5f:3H2;cOF.bf0f.W(\Q\Df+4IF-8
OJ?N>N:FYBgHBM[F,c^BVcVe6D=#0E]eLab;7)eVQ[V0>/&WIcN??),edIdIF3LW
T=>I7FOBI6CR[fP40FVL6+]F&)ZKKYQK64)gWTK/P+G,2@<-6HQ6)V3bS\\+GE+5
gN^WLcRA,M@B(8O5,#7@f^M9.CS4XQW^P0Q9HXAfd(?R.[8)IF>Ob+6)IV76=T@^
5X^X2Y,Pf-GB::e,,[PE+95e?YC\GTGe?WMXT<0\01,1C=+@XD[>QgB4LOa\33?J
Y,3).8M^gLUG.Zg41K;OH5cY0H&DV\PQeZ@=1+X])2dWD:K_ITW.\f/N154[#5&O
1GfT?/>+I>1E,NC_\+E&;UV8e2O/fWd+e]?b,)1UK6D1YgOANQW1bQ.J_(>;1#XF
PATc#?<A#FW\[BbTF=LL>LFN53J>(cWV?M7R^PTY-S+fY2D_?SV+<CWBPQU+QD4A
;\-@\<Wa1&-Xf?VR]I6HX&=U/(I\4_;G#c4a12d;NaaJDRRD,1E/N5Q76.]KKMO>
YL+94A42O#c9DVa/g41Cg(e\FEUcLb2-2T[WBgY76^GD]Xg7f]9:1-P&?[XH(VFI
X8F8G0G]EPN@OSfB^T1P(14@>]/O\T>1HF4BLGOe&T1cTZ]K35&U.:gc_e(/^-V@
daVNgT\BRX&aJ5WV+cCG6#/FD41cHd2XCTbTEC4fdc[\A0;Gc57Kb91-)1ZYQ_8A
H>XIU.e+Q@Me@2QEf4a?^JbD.(RLE]dK05_)8W^/eQO;Z7D_[L\QC2+PSKD_g+T^
G/?(^1]OM?U.&3C2N5X8Hd_@7Qb[JWBJ;=A^XG.eYf,&DA;E1DIAAaYS_?bH.Z7d
/WV\;).V9ccg.a;E21gD7g/[c@9_7I&B;Y68Y)>.\LWL_)I0OAGd7ES_KZ^<dAVB
9PM7M71/(0b?B;gfL73\(PS,)gV;YIHY>g40_@XGbWU0RD=7OB=]e\#f_2_XBJDS
a^C5OY)EQ0N7?#aERRY8#T4273B1Ue,I^-aJ;X<VaeH#\IA&6@-GN&R7)4dB6[&4
.5J?0?L^F=_[8[,/85[7bE/SVQDceB=#F]I)gW[O&TF9-KXN;D>G8f^Jd6.747&4
7;L@O=CFZ9a-0P5gcKY75J_Q;W=6E6S0K2&\-GTXTVPXd9TTH6M,_<g5>G7=B)6Q
PN3FO]H+2f.1TJ(G4IA0/6M;aeK5>)S7]3d8]2@=ZD::^&#8J@4b5=\K3:aED>1,
R_P=SBM1R;W76+fY_60f3Cb/-4Cf,K2R@g?;E\R/NS(,VZF:_64?M)H:e,-Z,;#A
Y2P<#HH1d4Q/02-90Q005<O,[4L;9WB+\F5<T:2?#0>:@I:04=S2d)L;]EXUbI-c
gP+f[-HU7HXF8b25>W,1SIH5>E/<INVP/-#5>Z6FfYJHW0MHf(aZ_M[K484K=MaB
,I;]A4X];f7ZJaaH+;JQ54&^^+<([+CO,>U]:>EdgX&Z4]NOOO,g41,VcYOUM4#.
-cKUZc2:RT=#=N_=4(.\Rb&?8K4a<]WW#\>(;@V]6^EL8^c307HP2V&f,@;/XPUC
9HX[VM/gg+9f,1P<QX.@S@#U7PN&J0>Hg6^UQ,aA++e)SVOE0W[5O.7N_E21J7+T
6#Z>#L:59\T+)3B^].M>B6LIa@?)]Y06JM,T0+,@Yfb)?05?X@Y7e48QgDS33[c?
=4Z(P<HT^->DRb\?4^2-A.WR&W#+FMCB?cTNO\9E,Y:,(Aa>@EXK)/3aT\eUa#f?
#[QA7ZRfWB_)LB4XVUNJ;U3HTe@f?Z8(V)4J0ZPQ)2M(Ya-\We1HLN@N7WKa.^EH
(&YBAFPf[+#T3&BL:X9gf#ZQ_],4cb615QZM\b,M1V1aMTgLYZ<\1+eBfU)O>Ja=
M]KDGfe.gHbOeXc:6[,]fLN<aSQ12V-7+.gG3MXI@Sdb@-29=M1O\8^)Ae]7X#\;
4X1WM&F24.V(&FI9TGI,^H,.-12Ee353.;=+VTY\=6g<gRNEP9;;Lg)ZN,_FTN1O
Z@]#,W@@04++T/M(K-/<;P-<M,UF1[;MQ;3Rc4]KX/BA/#@A:Z3<9QH>Q2fEc:7O
BSDPCJXHB0.-Q7ZN2A_f1#<bFV3Z5dJ2VF?,-+EcQ@[2D9,:Kc@[5fbQSH(6L6[V
cUb#UJOH+2>eJ8.eNK72c7E&?RaS#[4DW<-XIY_Y.RVAKH3;N32.57[/:GK-.),U
\,OX0&YM6baM;LD,gYb<\9YXJ@2?V;K@EH@WJK3<4O^<72@K0E1^cFe/TfXb&7T+
7gQ.e1&bc-<O>F6eeTF9&4ZP8aPAVFWA7:53.cV&<eAT0g:24VF4gGYZA,N\?YX8
@_0Mf(12P,7e5WND@DU[FHN.K]11gEW_ZM3gJ@J.dEZVeQ8T/a[.d/B=KCV6;fB&
LY7(3;=^72J;C#)1ZHM#=);Oe/KL6gV#R1660-\F>KN7.F#f=QG(\X02UQ&E&(ZB
<,;<Q78Le\BBf:Mg7\^6EJb4/a/(KU]/I8eEYK0g)^D10\R5A^Ia7b]#<#5\f9YR
29;[T6RG?/.&MHV^DE8B@EIZYUXQF-b:eK1aT-dA1FO:B3-aL@1?3BHMD#c0R<3&
Sc0R)?gABg#GeEU9SRMVE&32[H?<IG-WO/&bIL(3GaTdNB3bLLN],#)NG-9Q]<B_
f/TL&Kc=M6/3HV6;98EXe;D^+BcV&)H4A9@W8Rg6#(XN_<)\M..^N@J>FG_1CM:S
f3WXG.M(&5(8@4EPcMB([_QOU&JRI_L4R20VQX(V+Rcb41Q0<)WWE3S#F8VgE(^D
3X.<Ye3d94QZ9#U>[^TbGCGQ\&9;];+)_0)Z9,F?;+1SOKU;aLYZH[Ye,bGU@gNC
0U^&?9RN>-dR;6-ATRb:,FU9R8J/HT=?\F]40@XYK6POS3cEEXX2W0BLMJ5SI7>R
6SORJ.LMT63F)@[1dXYHLcQc\f^ba4-3<efP.f^#Wa73+-^Y#Nd-(f5eb+g6E[8a
KJ+#R<>c5JL+X\B>+Ua4I>3E7)GDa35?KYPY?7QV[R][HW[-2GI=0e@L35fWdX<?
JW,A@-,H3<(c@6WB[(^/[)EM(NCDJ^EMEN<14Da6))XG8dWeWA#?>SYcbb386)=/
J+,:K4;U5+e]U?\D>Y8<g^X/O17a[H5+dM<MZQ-f(7.,SCIU]5dfP]J=0dEY84#O
H9IRX6#Og2)A[1FKM@f[gKc>bG+2<Vb:]4,/K2VH7Q8Oe6XR9a,(HSd2]&W]aTTZ
aQF0_=VU>.7>=<]G;OCO;R>dM.9\;J_7>+=NYN/Ef)K.bGW,8K8OJ&^K]T5QdEG)
Tb&@9=UA]<?<T.@DeO0T0gbIf?0\;)9@D9-IW.X)>:9Yd&c].UX-E3PIU.R&]7/-
BGUeQ<<>[/32FXXLMS:@<Y(a2W/=>faO?4b.f[<6Q?[@Nb:K7Wg,9Y(baIJe=RQ(
\d2PcD(f5WZI82Y)Q4>2R=4Vd?#+Uc(QbgZ++13c-]^?<PASKc#X,[006d+I[,ZR
bgF4DDZB9>1[T=?;PC[DXYTL/.<4@Wed=(P3BYO(=:_L3d3Y=9K)b\-_g3Nda@?U
+;I9K#-M/]>-1(f:N6;5E7GWT?BRd)1JY&VRH32.4[CLQ)=2eC?A<V:M&:6V\6gC
Y[W_]ZCVNf_B/7Bd3)&AAW]cc&H\Qc9]_;,#UGU2I8TJgD+a77+ENA6:_<0_EGSZ
((\CZ)O,=Rd(9+=0:C]YX_aI@3QZc>.EAf5IdKNM^^b/=e<6?0ERf;)RRQ>-1&M7
LG?04,?)H89P3?NCBLV,\H#+6\7G,b:G:2>b5A+:T223c5W>HRY#bO=XA#;7R4:J
HBS\=X4//f=,IO88F.9Q#a<,FT/T;FL0V,F@.V1JVf[(0f0d)f^.K/F^0,X_;FeR
.QXd]#9S1bVWMDcN]NVSKYRU:_&CG+;#W2;UD#QJO=VJ/8ZOC0GPPNTPS+(H\(23
5+R0+XD,FR7QN::\[+F_4g9Y=5--D@&b8-+]d04XEEJ5Gf\ZCG\R?VdI]KR[C88K
9>-8ee-=H8?.C,;\DDLKA#OID2R>#@^_[,W92W#(>1f63\VD3YD-LBcO86V.0LUd
6:0_&/ZC;&@WT0J0J+EFQ2A[#USQ2W&K1@\M7M0ZGNW0&cR^7[)ESI;IOOW.-4b=
c/3_H<LQ]Y_Nc>I=U/T^\J;4?FEb9VAP]ZWQ<W90C)5GM8bcP-]^.+8ZZgI?=1O3
O)BE85HP74(39J?HCL-W035;Ad=1/;4IFFE/fK1-?Ig#_45XGc2?CEOT=VfM+g0R
8bC@&[\WM<T/d7ABMA_31E7VbOA1Z]AP)MMEEXEYZ61SPV^\AL]dF.AQP4(VDGB5
HfVZ#_,:HcCYHgd8J4HL1&c7d.IPGPT?dbb&].(3Mc_87</#.VXg4dN@?:bdB_;&
2/bZ[H#FHZc+B5W<<EGG][7N1MSd<da-/=aH:ZXda4:H]_EU+B+?G/d?)==SdX\E
+D>WXYb9VS4g#bJ83^>Rf:S#IV+IPJI/,Q=LI<dBS5RcH62_Za,,f58F^2NK=>#Z
9:E^IfD8F[D(A/DT;959.&(][8/#A;07MeGBUA-@_?ZgS-2D5Qe:9fE:9M:\IG\3
[cPd3(fd:H4]1O=PCG/Ee/S][26L>MMIJY]1eaZ=eF;0YOIAW;(JWMTgOJ?U6.ZY
?e&D0I^A?dLVb+>4PgOJON?GgJUZH3/&=W-FB@4@(UQSQCD5Z[IJWAI1;).cXT]M
7L+fgT2B&6]]+RbF(O=gIag9A3I(,1[C_B5=d0VNWb.==PSH^2\RU^33UGH:L5H?
SGI+.N2\N<2V=P2>0,B])7@XQWG_BYaK0_#\E<?7f?+O4,cO5(N+XV80L8:4_B;]
WNRP?EMJDgHFV\dZ7Dd7(V6&(0LAT0Va/LOf>dL=S@bfP_ULg:GITg-.TFM01?=d
6gCD:MVM(([8+_VfBR+KCS.&TZ>5EYAPWcL,TH37I6_L4QPYKV=eX/Y7K3R7]\d6
S]c@X4Ec?FHL@#AC@<V66P68d.f;IB]9f3;LTL)P3ZBMR1RH1D7@_U<IGPX0=UcL
2da3R3Q6)?VE=TIC?g\Re7L+OKR\dD.MBdI#3,AS@:U]9T9SO1BHgGf@_Z?6BT4Q
LVL)f&W@J(Z.8M/&BHHP:b=A#X5E@=WfMcZ0GBVX9[>_D6C^B(JFV(S&Q?XD3X.I
P:6W(e+UP(>0XfM>OF13SgU:[SJ@>7NZLa9DcY,Sg4QI;G_)cJ/\T(Q:ReOVUU0J
CW@5DUGJQ)ZbGDX7<7OMT47be8^=[:&bS@M2]YON04^&68V-F?=G(F>C@>WDRP2&
FP^(N:29XR7@/O[fO^ETIYM\:ZHBUDAL:_F0bH9OFa)?deW/=g;-QGbU)&c(?JA,
L0-D23b:9B;Z],)=&2>.bUDP3aL@AMA]IUfdb65;U+<,K35(g8gR_eIMY0N/R^EA
dRN<C;EeS9aeZHUM(U98<LW<0=:,_,IP=ZTgRP>IMYXZ9)beYH<RH/dfc#W;PS+]
KQV,XUB+9?)LW@O.bY^U&N#N4F\20K:TOaE&;RIYN#d,KHG(^03<74Y[>TUEGNC)
4cR:WYQ)(5MX9NX=10,M0e>&7OOLRP/Zaa<._F,?<Qc#=8Cg:YJ7TFXK7aQCGJ.c
GK]#?SMdN?/G=MN>NZW>G,#E@cL4b.>&J&P)\K/c]F_47>8-KUZZ6H#VB3>;7Beb
OgMP5UGBbM5D&=gDO-e:Ca2#g/cMD<GV8TX?V[+(741685,Q4HL^KR9AZQ1bSFQW
MX83\[86_7^;-)F?4?@(Y6ccV61(bB;#CObJFWI7/SKNZ2eA&2:[S^PfC59>EXRb
>>L/E^&<TSbA3]1CNLL/[ENH>C,G1HU570HbCTVQgP@4dc,NcBV>??M1-H><b/U]
W0HXM;,NU8N3aCX,BVA@d8)VJ<3P>#gaC:QgIMJ42Q,AI]-2_30P7Je-eE(-@JS(
Q-?9A[#&4BVY:J;b_O#B8<+ZHHc2KT98B/8)U>TGUQ66O8:Y>91A>+42)H/dNQ?=
9c7QFLBK#+@L8dCEb,0NN7=:D.g@P6_H_X^Q]2PZ//;Vc^&=LTIL9+aNP,JVa1-<
F(&8/bGKfA#M2H=+4T2<+a^6,&;<e5EJb/EE+4LCF0G@B)&O<JP+SMdQZ(ZK?B8?
>5&;a+\_eD_d#JM=?dIE@ZS;<-_/8#GDDX4Z>e4B4.INdV#&-F]DDU)dXP4cUD-5
0>AQL8AD92O8UOa0V[c.5?82S0g\e<&AQ6@5>D(FOY3&.JMb/.)F.aMcB(#FP#?P
/&9AE)d?=AI4I[Z<W_dP>]WA#-eU&G/J7^G3NF4-V0dQ0?2cSEF\(Y(KVKf2TY[0
(=7AMV61Ha9/VW@fb0Q)3+.bWV+WX.X@<(5Z;NV>IF74V<eU[;;c,L)G\W_CD2Vg
](aAe>dB>O\-/\:Da#=g/9,PW\=-BBHXNJ.Q8HZ>B7J\=[?DB8Jc)2TLAMMIUL78
<Tfg[40a65,)/A@^aSTdR]d_/2.T#?JCGg)>A.E)d)5[gTf((Eb+@W/CJ^O)W/5O
R=cEag/SJ6PNb;@BJOM[+bI]9I,Y&6?YZM)@dSd6b>2F0L7a\CN98O#QV<EFM9@3
Y\R7WAY&OG^K(H7_6]STLN,ZP/WA=?U\/-S_O01b3TN@J_B+?NBOH7\ANVG0N6O5
dJ]DYY(7D(H3_^M2eEgICO6[QE2S9eCR0628ZVOCWD2+MDY=;(:b0bc_5f1S10+2
2O8#+4>\/M/-6eT2YFd&5C7IQ;X[@L&KKfe))4Q)YJ@fb0:A;e6-J[EI4ABYU_cd
DZLWZMLIFJ1&0^P?ccf4JcAY2AXAQMaLM<b7O=NS0cTHe)U]PXOZ7/+cc_)=Q\MQ
G0],eA\HW=1C>N]4gWMT4\[O0HO_7SY,8\;42OgO:94Q[KH7K;@cQK#A\J6&A&VT
+JLI-AI1E3/BZ=?d.P44+X[Q/9A73>eX6T\8@9T)G)FHTc3agUA1AC[bS3CQ^0P9
Z>C#dR;Ba_eX;MSKKU#FcaJbf2Q5+:^&(dK&-A+1O@E84GUR@MPO\gC>-9Ug.Y5#
fP?/9+M1YKGC[<E[9ZK+QF^/T<5gVMQcPd[We)<,OZL7H_;39(.NKcJUI7HG]&7X
<73-(_g7A<7CB,GE#ZY_3D(^cY.C0#-9)Y1QPOXGb,\/Y9C88b,U4g>Z-6VDCMeP
J,-),TUSDP;.gDE+G04;Od5+9=DVT;2c.Hg)O>/a_8:&576&;,+D<7Re0AG(G,S\
7IcS7G\#&>M:e=>MBP:;R@;0P6<_gLF?0<3G:5VAFO6CJ\+.X68@X+@2fTR;NQRV
PfgY]A[X)U.Ie^)0dcKI+acTG3<,XZ^Y?+L?ec(-T_-)3/UD7M&;@W-ZCW33-</4
KW9_\g#g8X-5@PY#2XBfQHRAQ2G(0TbPG@CA7Ia4->^.Z?<C74I&M18PWeK2GYB8
00IK,5g,#^/>eB4J>OCbWOcSfC_,]I_KE5a\+d#W[E\C7d5^IQe+6WQPGBU/[.SE
d<SQ.JL>]&=1Z[P9I@WQ&2-AC#UO;<g4O_6<RWUCb3aSY#IVb1K,?EO4=aHeEL8T
Z,O(E8S:\fb3fb287]71_fRH&57cWY34fD&4?,@YM^&Vc(8;VQ]N)ZeZ>e=:\Mg)
&EE?W3A.aSWXMJUEUG.^HQY^cOcE@,>X8-XMf1VA[PX5=+MVdN5@WKL,6?EZLD.f
W>3;g3c[A^2;I^B7SHG^a=Ea_\XOFY)9[N7SDC6.H>C,=Z)YW89;Z[RH[gP/N?(,
:[]DJ-:G;(B_4[+U-)9[)U18R_0V@4ZQT3K,+LI:b#:?47)M-C-SFP@VWM[VC^MQ
HN4_IXfB?M)UPE#)Q?4K3eRB<X=MVIACQd^+T4P]?VeY,1Z1?2P<-#e/W6Y#?\[Z
V+X.MF7[ID\PB8?J/g:<FGR=\:JH^eZ\CID&M7MW#ff(O8BTW#c]3a9VP_]T;OI#
K#<X+2NJYeS\I3cO?(VWdIeV>cf=F?ZRMYYLAa/-J)[S6;f&8I#[KOTc]6^e1:Pb
d)^E+Y[6G7/NXcBM7I6A]<)<fa)3N[dg];)Oc8Z)/30VFN3&2CGHPAK,8WEX#gMW
6aSWQTV-VCRH&#(0C?6Tf@#?61J6<))^#\OUeG&8)S6f)a+S[^aeN7cA4WPfVH>f
\36,>aRYC&cRK,2?&;BOK6E.3ZEEe#Pa.c7-&&\Lfb.7=:S_c,#_,W.::77^+X]5
Z_H=B,MbF&CDEMDBL4WY9<=FM.4a-I051c7EK_&&YaCT&/N5H+DAUF1:^/R72@c(
S8T^#.:1)HHXRRMJ_#fB,W(ROXB9MbS<UE+?KfI?&WMK#5(G&C1Y&Q;NJBQa;60U
)Q@NY.X?\C\GRG>NQJ3MMO6KVU?9[=8O\>>?+EG[JC0B,D+d8d^g+eV(Nf;4+-Z#
4E(aX17#dW+.@CNV&IUN\7LE+RV<;UTWP/->(dJaQ^eB7JUD5F@#A-L31,6=)6J\
;b:1#<C6XA)_U;KQ<K;W;P?Og2dAcYWP)-J>e)GGd<cI)=T(PB(]9>;OY2]T[MbI
=D9bW6;BA5J^KaTE(ZfagDEM+[2]RT0MV56+IPG@8UP[/Mc(Z,D5UWDPMZBJGGgX
.E7Q:X>,&(68Y@IPZD[)/f::d#aHR4WD>IXM<V8KA,R3\7U+VQ=(.TUb2PBOXAC\
43Q8I1aI&e(MVB?MBDB5O>TGaOI5-e>DYV#g>J,8cGU=Y=K4K0/O7aPP2LL7&<fA
:9EI<=bKX:aOB^7#WY517#TM)Q(>Nf,^fX49^3YIVO7YU@:Ed9N68VcEJLO2L(bQ
=2M==bGc==ENa2b@YA,L&8[Se)C_CN2G(fB#-AYHf;/>/PXIG^]N=XNOUPES?;O-
UH:fIE9ZBa<;E^G?HJPQA4&<34a:+YYN<(36[;-I\0VJVQ>/7KQaa&[C8;HB,?8D
-f_;9NZ;4MME=;?RD@C5^PP:T7M5@1U5-g=FEO6Q>ADXE0V,^fITf9.Y>GH@GX9D
./8A#/U3B;,VPJ=DDRU5/37YO3.b(KL7:eNfWeV,CR-<R@Z(BG]=H&XTV,2+ebSR
FcIA,7UF8IeNU2_TJZ&<FYXEA&MI@&g/2FI+G1[eD:74Mf3e4]0;5J;U2bdIYfNK
98N;UZHfMWMF3HJ<6]5V96\[WAO^W\;QXbcKQBZI0A-T6DKI;O]^]?I=HTFePB^,
XJf=Q;:#[(M1\Waf#FQ.M,:@Q_M.^H(Je#>9_B^KN98?>BZCGd8(I8)a=3@7N.HQ
@B)#ceG1/XWBYMcS)Y<#Yg<bCJ5_:UX[YZdEd-d<F5cKX5)]R]OeK@:)Y&W;\U<^
\eIGYE^GA^ETIIX4RH#[S8R7MJ]d(Z089O/>fFKa83<L+]a8b6#NF76\TT:A24;B
3\08R:gJ=ZZT6Q;)OE@K=I\HYG@,>FT<a)Z5\[@Ed+^bcL=B>6.SeKX1GG:fUF),
(XAfe)0(A64GVC33P(Q[U8-Q\+H0LeBf\cC29@5ZKP-Lab]LT+8J]#?41A3XJ7N/
<UX=:WZf+#-Y#A6XfS18A/I(#QKcP,bS/Af./NASKBENX<9>UNURUNb]9V@)Zc<Y
-@AAGL6F-(SNZ^TK3cS-a=LFQ_D60bS8;IT#)&Hc:U6@1AUbf\7e>(?7YCbU6/NL
A[OH_4N#9L46&^ZaGBM\\4K;:6?4>[,c4Y+fC#.SP]E_a1<LQe;ODVX1BQQ73>fF
-c,<L)dFMU^7HYcg4TU;b<M[^RSX]?>WXKOQS63?]@K=&=&2;FaLCbL];;H4-S#N
SIX8+aWHJV(+;,T(f>b\11^^H7K(5+AT5/]5<V)(Y[:]1g,BCG.F)YHfTdND[\+_
][K#(M;)MR(a/PP=TSg5Xb-TA,[1.Fce[Bg@+T:gTC.)_7dU6/GP5R(e;[/S:^BH
a5->];-YCNK=6]R:V8,]MK(;+G5H#GY2YNYHC]>MC8;^Q>(-.AeFD,D>WU6Z@<R&
[<b6G2W\8R;c_<+SQJ#Y_3)Ne\UV9Hc\bC=[E+9+,GB<GfbQ/9cJ&BF;D>@_90U\
,aO[7:(8Ag^(1;9Q[,;<?K-eOH[)20G@=89+O>1KQIPA>=2YS.V[&T)a4C[D5:UT
H7e.;5-&YHO9@CP7UWIY<UN=/80FQ3Ief,Z5Z([Ea>GM/<O)JcOfO0)?#QE;XT^U
ZMJ;B1),2[;>f14-aKb?NWS=9/MZ))d?]:H81,9F[(BXM=)M\7V\c\dP,SPa?I&0
.g503cZ1J.6-Q1@<_,Q,IF/\ZJ^g?BdG>2bK50+b#A1M<]KIc/,&c1#4IC0_^dEH
c\V.#IX&3\C>[1H>_AUW3dZ+ZQ5CHZ#RX/PV03UM0=Wa<898P;^B4d#K-H<@J=6[
Kc6(?5&QYCA_92c(CKDN_\5W(V.IeQfTQ(]_7EM:T#IZ#V<E?C;gN+\EBRDZ+T)L
5>egVECL/J&g870ceef]),<EMNM6GDTSBU95TS2b\S6=:.eUb+#-W4B[CMAZ_\JG
7>K>cJ=ZY_@4UT:Jc+#A<]5:ad.4YDaVAOMg]3e-2397F+6WX&+KgL/P+-]QN3C?
EL-9<1K3?7CDB\20[I3Nc_IT4FK;0,&0A-80D8aW99b3=3bI_,M3AS@f;\[OQ-I-
OP?;V6;V:5[NWO,,=7.)0d?E>]9@gJCgG7d1AJQ0Y2<=\BWK:U>]?67FW5:ZVZGJ
&GEg\Od@I\a/UH)&bfXUXa^PIW2,(]bP+JHO0DKLN2cD2J-/B#ZG>\=XAc2KC#5a
P,X\,ObMZ>SVC@&B1J5dEVTbZaNaIU.)YGFcVX#P)^UX#92W=(D^J?2e1^X;ed:]
,QW=.e2\_Yd@.#FME7>NJ2/N/R,5XQN00f1=Ab^_NW^Y=0T,<_]a+VWT-S&9)T0R
,]-TaA^2H9=;.Gg^9C:Je3^QQI^f(E7Ib2@[b7H:TY>EPE]Ka0E5dY/-B]KaY.fD
M7#<5(RagPE_TfRcd>TG#C33DS?Lg\YFd?M8B(_E9K&2a2[+P6;f0L;=@I(bPK0J
9b[/N_#8=1R4>WPSA83(eE/(\U,&6aJTM@L?&N.a4fU/6FeMf[0FCM<V[Y#f4)(c
a7J&bL1a572-9AL^]>PLW\;8B2^YSeOW7Og0GCL@O3eOgR##CCO]-ZXPc98@^]-9
A#dHb0#:Cd=7ZPfg(JB]@;&eBILBM_dO=H\EK+N;3=R+L51EL7OaP],LI^)8<1@R
)@FDOf]6K;YTLKWc;:U]NdL7d4dX)7cQ))DRfA?^JgXZA7YV^VQJBYd\Xc)aHe&0
0FBdf?+)\JMOF+L_]Fgd2J+Rcg47?JHd@3eR@5&NaL5/)0GM(,fQWTOc7]ga(3cX
2R-_<2Mee8GNge<Q[UB/]\)W=F#c5^EMR5AEPTRR?]R5JL7-/5#Of-8AK#E0XD>T
+^_&bOOOMWR\4NS&28T3_)&4=GLf0-CA._.6VJPAC;6cD]CI8#OY2f-Z:febIPV7
\PF=@P-/=WZ9&CTa+ZX#1)/NJ=I912]OaLX&H]V6MY<QBKI1KOAe()[[OD@CLWC9
6aXFSKY.2UN2JL#_G.N\(Kb4\Z@[O8,NJ6dTGOEfYf]E3Ib=_cOa5S4][&X<Qe,_
b?X.5RE/a7V-H9DQ]QJ1(FFc2V,dDDI#].;F,1Z\/H_dBD.Z#&+Rb4Zc1P0;A?,S
X+U6@UgO?#)#Q[[a1NCY)GFeA^4(+&L[[2T1<JWgNA_7[Rc&9IQfL7,T#GKXUQfP
QO0:,NfN_eg<TRZ0aeV#?0+HP/f:FfHRc/?;-+fDX@S#3eR]g0)H+b&,P];Y&-(F
X?e&OUPagG[P):O6]80WA+CdSGRG9#BX&8=.56=GD)1FFU4^C5(QH20.bM#N>]O4
5PG8;R]+XLG550(bCKSRM&BHgNAP9ITN/\Jc[A6N?Q];;WHb<W0E5\dL=2E^&^[)
[/<BMB+\=6O)2.6U,9@2Y,0J2O/2NH=Ka<]B,g.0S]e/-8N9E&XHgQ]63PcUVG0&
-[^3_TI#UcAM;@AdE;WK<YP^Q.9YAd+dG7]#]I,(&S@fYMTWEQ<FBI@)M8gP,:<G
IVFB5MQ7IADB#VcVCYA[T5,R]C2eRJL48ZUE,eRJ[T?&BD([;d205,3LU&9WRV<#
ODbL#[</;O]N3P/)&B9KHYYH,JZ2W3F</N@95A=9+>f=<:>H<#0bZ28+QcD-X[Be
d[IUM6:Oc61[_7MS7Q-b0gLXT@-W#/^A\FEgUII8:e-dH^4P6DXXEW0[L?A-9,cJ
RIb(3#2B2141]_H^&dfO2Bc[<2\Wf/M^0><&LTI@[NOd&K_[2gN?LYVYQcN7N[=Z
c@(?feW09_]gPV?CCQSQB2T[7Je#20PDON\4feV&NW<,S(.=[+^3P947K(\Vc(UA
EY@aeJ,M08^4X/BE>)S+YP)6HI^+Y_b>J_Wc:PSRa/HV^ce?(82FP82e;4NZCFL&
TW0+KL+SD8>@;J<F/UQF_^X])E[@NgXJC<C-07a6/^AVGYYJ>/dQ:0Z<YNT-9&Z>
Q7)_;>Z8Tac8<U5M?1RN.Bg=W7We2)S,?baGT@G+dFB[[&JVI,6AU>eI(ge3>0N3
:@#BJ+\d3_-\YMd8Y?ZJ)2-RA)c(&A#IZF@@NE<-:6R^@E=FIKHOQ.G1=@FT.0Sa
#@e(bL[:,FN0SJ/b5eYbG?5-3&M1MQbHFE:dTT0Y=5+Q<;+C.=g(5,>VcBaOb<NO
ZKG-C.<T[EV&(EI(#XNDdD4b3fJVHR+Re6R(UY<,e-FfeUE56b[=\4SI:CTLHA_L
3OaY_dX+I86^0c)M)][^R)@>T#W?fB#W^,cW)DNbca?@E(2)VRT+e;83gbWQCH>M
,H)b&0<11\W:8.<ZCLD]gYWA?>&DCXF)CKf#0IN48-LK>1U,7=P_79F4?^[]),e[
NTb5/E0e#Y0EF?KUZAFeM0I3[P6UZb?.3DIM2eZ_/TZTFcG^-&Rf8L(S@+68O-7T
26/#/>Z;J4_3PCCT)bW:fO1?[bbUL&;3/@.<T1G_Rg=f5#E>OU#B@MO:49SC:1<3
BSL[0VgT,-dWU0YAX7;7/:Z:_H]Q_Z[:?2<S@dYO@=8\DN_e58](4_7V+;>52J9)
QPV[XFY83c]8(4>3]+bYF^Y9[N81MP2L]@9@;Z:7[ML^U<I#<U1MTU\K]9^bSdO(
dAT09#3E5CL.]<_K]+34d,5R>\^XMW7-_;\g9dQXU.G[.]30+++L&F;^0JPW8_d&
Ob=HIA;ec<+XcIH9U,6[Tf?(,?Ve2T3gEK=a-AM@1OeAN[E;S@)d]L39b=1,RA[S
AeNEB/D#b6J67,P9:-Uc2M;eaed/8ZHCG=^@\E9La0e&K1+#9;A?MT=Q(C?.aJ(G
3;&]=W1K_F?.J_RY:DUL=<]<3&bWgOG[(&RR@NeH[XB8f;:4FZgJVa.?RDX4DUdF
7)ccd38gL#J&J=NReP5E231;@7#3@FU/O-LI0ZDfU0?)3SeMfH3/J/X,NZ-55gQD
2aTW/bSaB;LY67K8CSgYY-996:&,@X>c7.E.1EJ,?/9V?Aeg=(@H)2;=3T[>S]ad
:1Re0(:O;6S5I,T<V@JSaTMY>aRQ1F\)H@2#8AdM-c2[N)Eg+1UA#A>/OT1b?7[Q
/XN8R^PSI0:F=A-S\HTPbQ_bfRI0M-aZ4b7M95U.H\-2@(1eS^55I+;E_dBZXG+>
>BE,HV0/dQ5eO52N.G.44\a,+A=/a6d5C]U,;+a5g4C[3TGTZeOCIZRUP_GAYQD&
;LFZR2@a[PeB4X6?:\V6B5&Z&7OBVA&_PQYZHKTfgX(3Y5Ze\2>Ag;0H,T=84g3R
B5M,5e30;=?:>BUg,VWMA8=e[[EYQYWIE#+]QFgT/U)+8PH]SL06gRS<YCfeETH,
K>N;#(5B1I@B5-UG,\c-+0:/<H=ZJ;&VTWgN;1B4;b:68eMJ(Lb.U6JWG:SgFL0@
KP25GY<&Zee]dQ#11#^_-=_8OJ:7#JZTY,=C=dSYAe:K.TfP0AIZ+a0OfC59NIBL
#3&K_EG(TFeLA4_8&d/]gZRUG]IPAW9B6OVPfeCLG60M79\c?[fL>/DPSIB7DH_T
TLe7NVN4:2(TUAM\L=>&0b0/YQZPU5g_.0B&607Pg<<H6Q<L\I[<(d7Z54;g)TG1
gJ..>F_SSG.f>gS--]W79A+9,](=aT:+=XUYG[3?<aHN:Y2CE^6S.SJ0d#1-T>:O
g@<9,U=#,.CG+geX9)6KAE37HPW&TR:eP[RG,CV+69\]Z,g)4C6>OR1K+9(:QAN-
^4gb]:(QTf]-.^53(\dSWV9Cf\3O+.J;\(:Z])RL)aN+f&D?(4V7J#HU<(<L]AS;
W22IdMH>G7F/+/-RWYM;@)Z0H4G,^F-@?cA^YY.B0EO7^LMQE?CDULZ1?0(L36JE
G;I@KJK9UEYURBX,BHSR6P&=0ATNI41?:D8P=Od26C5.KCFM(@#7/1fG>;V4ON4T
4&H_5GCT3#<N,B;#.TUP=5(&B<VdJ<fQb]C(<R2f9QY[_-+)85AU.f.2C=\-WM=J
AGY5_(Za:@d64a?]M99Z10c9\,W<?#:;<ZE(=]X64LU#=/@S\?ID.46P10I5RT2\
>eIZCa2cMF>@fK;cgf&5b_48N3P#)5Xdg=Bd(^26S:9b=Y7H?_>c.A<)6ST+M1?7
[3WS1b,5@==c]U(9Rb_RQ@U)4M(HbfE_9\>8aW894,82^-F7B5,C2Q2Tg82TV&Zf
Y=_g(aT\C7/C:\A.99Ua:W9\]1g6:d?QH>Y(S]bY#/M2^(gB[<c^[WUaRN#eDW4P
YebG=dL#?YaOb]\L_)=DUCF46[Cb]K(@Bb\R9dK4/@3a<0BH/1fL[=UGU[F3-MBB
Iga+fY,(@)E/3R>1R&aJGMY7a(bQYf,[NE]\+]R8g7]/7WNY>E,BQ:O[1IPFO9PV
4P?7QY<=;3\6Y6X2KIJYbbT@39/14@,8/F>94g#Cc@GE5HHIT_SUScIV#JGZbXQ?
&e.H2dZW6K@P=EJ?+AJ6G\R847.QW&[NK8Y+e4,;(N5WP#]^F2Z7T#]e^@?5FR[D
H>V61V[__N5UDL,JIDZU/Q<dVL@SD=VHNI+3+_ebZ(/4B?a/+/A[BJBGK:=8F:HB
J&J[7A3aXOeP,b+ZU6a7W8(YJ\JGO,dAbZdDQK:Z0#E-X=HccJ>.Y3KNJeEe74;:
FH?KJ:F.-NTXGEg&(-PH<:c3e)dc27+81G,J,J9+553SNCdM_&@IS?TV(T#^D^9@
Y)bGeA,;^-@+3>J_8g2^8aZJ2:^+<U4.cSJZd_^T9U(#1e-;c[ANN&>[L/:@1I.H
I:FLSQbW)/c4,Y4/db2Y7)Fa-=ZO5-db]<f3L1G##SAgWU(9&gebb_3(@9HC)YgY
Z\KQ#)[2>=?Mc=#7AP4+Maa&BfS.>[S;F.fdPU)^LJ=\P6:44;RCDf3710G2]G9R
GPDd/(9.cMU-c0A_NW]91@WM9:^8(&YQC0W2;b-_,J0X#]4JX+M@101;Z=8>g,aa
NGQ-cJG7U]9BE8@XK1HQ+;J:3KeB0JI\IQ5_]U=:X3#(Q1(T.P^gFUaT4B50g5bF
_7SQ1gPW.e4<I+;.Iaf-QJbg&5MDR9#]UU\@-[(]JYdWWC#LdTS>VbEKbQL4L,MG
LW)K5LH8C0H_A=cWP4g75Q9c=a6Nf2&6H2WO6]K[0MV_b)UcQVEVRR-<;]>(6Q\W
c@T3<^(),Gb?8>G5b7e31Nc>7;^\&Cg?NB]AXAdQ7Y2>CeO#CFCB.HU5._=bA<)F
DR?EJ.&g)7(50?@XR2NdTDZAIf]g,dM&@7SeFVBU>F8A_H.R6@WDY..5P37S5aQ/
cUaIM:ZceLWe),g.;#()3:U6W[WZ;5U]_L2F2\,2aS.]:([RP1H#/PY0Q1fcIUL>
6Z0(2QG>278&=4(EEE=c8EX\>495?SCe+0QVcP0H;)7N(dBe<T-(ZJ_S&=d?G7Q=
81TB+Bf]2G8P_1fF^/.5_UWB=PHgRNe=,e=5I>/L<EN2L<UW&?YPI)Q:M5/0=IY0
a,c;;VaHNS#,P#WY6f\J@W>(>MP?(5g-[Ccb0]DJBX68IC^]<La.P@Pb.E?_AcVD
g6g;(bY_d1B6fF2Z-96#NEKD^:CI9:c@D(YE.a.M5:-FBWOVO6X0g2E#(H1a>#eK
N:5M2=W83D)9&E,BbNTD:^M.f1KV29AIbV@[JXNGc;FO,F/#WVB1A-cQKW+._KRQ
V?KF9d2:DVH3SX;+g_.d-&)<)BUIGdG=bG-2;(SR^):N5^T8?G[6EH]ETPX=T@2f
?A.H-)fBMTdCYRVg4A\C<,(fJ)2fBeC0TU@TaD@H#IeQFEJ7YHSbV3C57;OAEASL
4_G/J#M&SV:B23M)^UHHU^9D_SCB_PKd)<?@Ta@2_T1Mg>,U)L7g,DI[I-?/(9<Z
4HWNFM<C.7KY&bDU8g-,Y+6.&_;/=0&.GG4d#IV<JVDU8,H)gf8I_;>P@E9IGd.L
bOBg?LRMTXP_6(J7A-=g@4+eR7G-SB@64_V6\:R4@X3^X0W.C<\@,4cMEfDN-6/N
&d(VZEM)AUJ@Hf2-BSXC\C.I&G<>5Q;JdUSQFUT=(5HT/<FfV9CZV++AHV=SHBD,
7f9L@LLDdS;WTY;E;\MNB\(QZ:dPZ=.@D^-61,IC&+@8J#3,47#[R=4,95]L54gX
8EbHPJ5:(ON,KgV<33TK;@M2\_[U9XM.HIcGS>&e\J9\U?-,Y](TJA)>CJOR@BL^
\0TBHC&:4B5#SaWG32U],bA3(ZBW9=-6WN]/WZ<_Mb:K_2-,(\AF#8X-MC7_SI_2
I0a2\KHNI.7[_SdOEXY0f6(5(AH_aMFVGD.GDU;:DKRNJHFIcWUgT:FLIMW-COeP
D+\TE=g64H4_JC)X?1Nf)fg&R=&,aS_CdQP0UN/U=LdS\JGQdS#&^TI47(N7Z2AG
\6^[;7Yb^6X>eRT[SH:Ued\_7BW0&(A2MbLbN4.3Y7gT:\/KI/+[X>1LN4YNESX#
(;a@&HV+L>A9SXGe;<FH^:M\b&)b]S_#b##.<bJ0Og\F/\)EeRc3T[fLCSSR=:<F
;4J6L[gf[O-C18\,W2DU/U<:(:)&8RR&,W4Z6K<6RD->c;U&M)]O]FcJ[91EJ@g(
]963901=Z6[9?]A5[AMCX.S\P&#<);H;O?U3?V4)-G^O9838&UA2#PP^>O1Z+&GT
WYC)1OD33K<A0N5X4;fC0WD<3GGgR->(:_<&)U8H/?cA/;R@F^a7J3FJgObJ3I-0
XC;.H:J,PYXZ(SM.FOIH5]M+8QN3:N>\OY1eDd]RUbO5[J<fMZ3WY_C+4:C&aZT8
=/?@aa=^aeTDgG/:.R6,/+.S=LSZP,e-1C5aO;VSO(K<RU3Ba=4TVH1PHGW81J_U
ZJbH;]VOdU0O(U5&P3DM]][18cRB\4@LMI3WXR(d4VBE_IOV0M.S9?QFL+-/K>a>
Z3?+/2REd]/<9&E7;A[?8L)(;[->TK_NX,I9E+/d8>MB?6=0<[(OG-55P5W;6\25
>TCb/QVf8YB?f[/6QbbK,\?2-YPb(bNacC5]G,P4IE7Q@67O-W+)=@(BL0PZG;,V
Ze9^S7XM>WfXSXb<24]EB.;(dR/UA[+ETN]gG\=\026e-1(0,E(-a;e,5:>>7Fd>
M/--J=);HLL]b]gJe3KB4BT/(bW<D2R0];g,V[B0bC=V8g[J4#1QEJX\;_B)D(,2
<DH4\NBX<7F)K5ONb]+2I[[,+g]K)XJM.P<8F4,26\ES.KL09LX=B^7P[OS@FR1N
\6>fP<A]GP6[69;7SU;X=d,2U0:E4?P,A\M;3^@XINE<8bTAZ>e3),eU90D[TE1<
:2c^:4b]:T&LKd/@_MJb_5,@76\gL]?34W5S\8.7++b)IYYDTN>#OJ.:35IEK]:_
2;c0YBR#0O]C=AD[8fDWW6B^:^?<8Re61Z^G@DUXLTf8J+U>_,e/P\CP=3-Udb<e
DWK\38+7f7eCQNT8HggHBZ^DQH6.9>=_J7SA6-Re&I6&L.&\S0=+X&;#WA:TaeHe
EO=823^gMOOONb;_F?R\@a<66(d/UQ)@51V:>7<=f9[R.Y;LL2SS.]X#)dbQ5a(P
S4DK:.T;6H;3+@0G(>TUF&0.EGD9MFO?>2ggOZT;1J-e9HVI62JQ.6Df#bPW,F:H
/)R@+g6)DR&S3]5PK2JN+Q6\X].E#8+:/ZVIJ</^^KFZI2Q_^2G[Z+H\a:5A1c^]
a5A-Q=I]\X\#]I<=^LB2W>H@ad,GS-A>?+#IJH.b3fU]=\B2\Caa?<5@9B/2aS_@
eYYVH@S;&5aHDHG0#M;,e-8GOc.W,E<0=XF7?&(g>TNda?I[\C:WVI=Y@^+J80d9
9-]V/647e+FP/OV0P\]Z<.e0/L_;)V.AU#f:9^Ra<f+H\&F+3g8]cTYJ8/]Ud/Y<
fMQ?53BV](f1W,OC5J)3&G;EN_3&RN1F9(UFbf=,@7RU?]:Nb+2:f(T)/WPfG0aX
,cDCZ&L+)bS]F<V)6SY(8UQ8Ib2<1PF8H/8gR2)59-Q^#Y3N)\Q^WW=HB/Q256:f
X.,QIU80-OJ+Vb:02Y::_cb_,WQDa8998,Q11fcR2+W7QVTg16E:87GU4;2A^,d&
RSP-,L#7aP1Pc+_25FLB+XEJXA3EP]=FN6WKQ\)8E[gJc>\<HJD>g<?E@&OS&7[)
AJE:9&.b&?HUYHZ&^-)T2f+YYd-0B5E.WbV4ROQ>g=K]adTaFSI+DM\feK]JI[-&
VBO#2MS,LF1.-b@OG&\_7N/6aEaf-e3ZGg95[O\N3][./W6]HCO0=T;A@R)^]/d=
6-XbUeJJWSe0RA>0ON\\G/7KVRUXCbK+f=6b6^8Ua&PP2]JU1.fM^22\TPMdDJ1B
TY7PDZY:?O,^.&CaO=fP.eL7VQKN=760@E#T:b7+T7.2dPNBbg;E.27\IJWC9g6e
K@<_#b<WGeLXT#1:7+-dYO0QYBR1[7UX@]Jf:5Vg=._R&S]OHGRb_6ZKUgD<KbUg
&.R5WC]\bE+e)M>=fCI7Uc[Q;dY8J;NBfQ5G.R9.76Yg:@D2Yd(MR_;51a9EI?CO
)H2N30,H>7W8daA]HM<S+)dY?@>bW<UWY0CV].)W5^>I?B]3[F,aA=:)g+IFC8bC
U)c>K8gf6@PDSQ]58KaV?I--ZMD->dW[L)@(+O_3Ob7NYUQGXSA4ZJ@7Y+7eD#AA
F=dbb^Z7[&D;,ca@Za[XafT)[K_I\\HWca;:(VYK\APN,;8X>.Z6b2e20W..R<4K
2KGCJW@Re0?J;CbV3?\/8?6>=-+IX.9@S^HN:dEA]PS2W?S20/(B7T;,NL4/D323
]>(POY9-N5/I#N,V:RIM7ROFCL&X.0G-caS3N]4ZZ0XWEfU55)8YWC_.E7+1:SY9
1fDCJc5N9YU8UCNe4G-&ZE.9W,>2Se?8S@?<-ZP23d;#fWdE8b6fcTa;:0f#3?N<
?#\,4CHB70b-G,/V2bGfGOH_g#I,,@4VSX<4LNU[)c;CIC9CAGSZa;Sf:bCW:DWZ
/NW]+X?1dgcNZaWW=P>JFeCTH8UT-U@HLg=B;#1W=N,4#WYOSc0VRPDN#Y[R7:[+
V1W?0A^LZ-IH?HEJ7Ff9)JID+gf4;?,#f5cYTIIAC<SCU&(1X.e#<6c,]XfD,P#?
N8XP;1_J/--588S.:KI@3[a1O\RN,:88IQA61[b(076<7;F\cC)P\&W^CbH7V[ZC
T@4+P,9R2Ag86IUVb_C?F=_#X^6^5AOXM#EZ@,-;gCgK-]6MOS.0ST8_AJ-E0XR/
dQ@\UQ=PaRY;9:2gA61(37B#<)5PZ9BI:\[FSCW#>CHJQXgdR9N2)_+Hc@K64H,7
X.F+Y0<;N4:&&:4O&20;E8_e-N8952RUN/f1H3HV=#FNT2Q))fW-&=Hd_:W\ZgTd
S7/Ae[A0C:f-b5S#J2,6<a?_Q@&^G;[VF1G1V6Z:6NU50M8&[7FFZGL\9gQAc/dF
a6H^ga8<3F:W5JS<-EE4C-P^BS_eZN,R2a@O3H??Cg50aBA57Se;e:<=]Y]8/_>Z
bd#?U35.BcL418EE5@>0:O74,GW3e._^8d09cQ/9FU5fDL.0<&dd_JMQH6c:WZS:
Q39a<TFZ8&U[E=QP]E;(Q1b;J25e^,WT5)L0P99)VLWS[>e_,?EVH]dPDO^2V&8g
2RU#KK2PE0/8+81Se\dL>>3M2>(1?O-84c5FOK#N2UcU/>5JKU2L+AcI[RO<R,^>
-fa&MVH<8RGNaNdeWa_gZRYO.2)&f6W67^#\/=MFb;:4HP1I6\WS1@U8>0d69^,O
B7IK&PXFfJRRQNb\fC:fR(O&38<a9):W95(M7Ld^8LJbBfg,MWI,IX]FdPU;XAdI
:_Y<b1L:[WDYD]ea8ZS/+0/<RCAT+>]>_YEO_@<>1JCU=2B2eX(NaVgO+UO,B.C>
R/_ZL8d9,e&C=U#c8Ccf;<4KCC>ECfXWD(-#@T#eE88&eQH=e1AE;6H]6T=EQK15
?DgL=_acB\e4&+gA+]GEf0:a6&V31KE:IQ4K+BC8:bC)I2dG<N.6>5=+6g,Fe>6O
db,X6N#S=T;4CW_[ON2VU]:Q;9669\/EGZX>6CO[N?PJX=_<Q@N.._1G,MBH@&U4
R,C/(9\7C/(&V;L-_1S,J7@#V;5BQ<6ebHO,dN;:FA?]T:6;8]BU_^_+86)>ga,,
>R6fU+X2N=P]-BYL/CTXP238Ed.)16?1GDZRaAdBK+AT<BO,c+Q+]=J9e2?D+PRG
Ld&19^ILHAJKQFVbM=EB16b>.)N[d_:Y#XP<Y,g\,C>J3LP<X,NXMF_5MKT2,Q5-
Bg(PA5_9dIH.8]U#1[7V)e]W0T(<A+U?be-<?1\Z]_LVJ39?_+8cD-&[IP0IGQ[6
GV[I@TBRU)3Kg+E-Ag^;8Y),D8@XH)X.T/gUEY,U4[fPVOW,[MG)L?TECEGVKF&,
^,B[CU4KAW@Q]H_:g4d7c&_=]&4Pb,QRe@INLYD/cfd+g_7GVA#5OQ80>VOCDC40
d;f7CUU5Yg1::XLHcUZAJYPWT#Q<S\J((R+P;1aE6cANXQ21?F5K[e9,R=\<9]bS
/F-]#e1<fK&gI]W-N#FNQgM@g3BdWL\L0a+fa5+JXd^+&F]P1X@aCQ3+=;^V6\MD
_;O>I4V]/BfE_S2Y#<eV=9[JRP1?>IH?\)Ne;/,(7R/DHTMS_T&M9[E@VVS-4]W-
Fg[T7=K23?2(ROO42^/HXE_,=5D0TT1L^<=CREAHM\MedSKIfK9g#@HZ7YIC&D8J
2JGT4Wbg38XE=@be.SQ@bD&@7DE=3C>ZRaaUI@-;Hag^XfB6TEI-3N\VW(c1FT0X
LLCb^ZJGW7FGY;ce]E@eJ0^(/@3e)B(>Z+L8?9QLFRH=(R(XX2SR#^<(d2-\;3J@
3?>Q9TU+e2)g^L.9G/WI_LM74\\UD_+^^O/IdKf0SET<;-B63Le.@0TO=a^#LZ;@
VAGE.2[CPWV>^D&5Xg2_&,<Xf;gBK8HT&Zfg]9=5Q98M8EcG9JVA6FE?OZTeSfDd
H]#(8.(/#CE6aRMZ7XgLfd&SH776d)./a-bN,Zb1\DXf9gBYQ-YG?Y_5M/D/d(>@
9W/WP03A#H;Xd]9+;H1WLQ>LHKAQC20>OD&D9I5d12\ZH_b528=1SJ,QZMW:4]I1
a]d#@[@[&F>9LRcRX?+Q=Q?-8J1F=VLN(:L#7W/&O2A;Vg3KB@1<g&@cdHF]J#:B
=]);T)^.:_L_VAK1MV/g68TH)Y^7UB7@8Z4cMc3f@@0VCU..-\LZ^d-/0\E/V=Ba
VQ14eLJ[?-S5Y#A80ZUOK)f<H^;[aaZ/GRSM;Od?M7Q@;J5[DG@EF&FJbDFEOgD&
g04XWc5Y&P9EJ\7N>C)AQ48#eC9LDA:>E>dGG,Y#9.8TaNQfHFN#:IDIPDMPD_(J
W)CbNR_[9:T<,_H6#@(0IeGDI+NBOQKG44eFGcdS(R/>O3f_\/e&(d3WW[:]12LZ
]D1X#_+C21CRK-TA9YggBb\GL7B;ZdF-eT#F^Wg/DN^1.:Z#9J9Ce>eBF_//[=CC
60:O3Q.RR<Ze5T^bb-YK:,5-M^<61dgR,^IBFBTBI\UHB,-62[6R0AEOO3:GMa]6
fJD)eK32XP9:;S6;Sfd-(1?c#Z]aTPc0\#40J#=?8:YO7e0Q^11\#Q,-,]b)c()]
7USL6_85.9Tg/\625-U3eYc]7<(M&WY1XV<f#8<0-S=c9#]L#>2YS_+L;Og<P&_Y
6bbAU8YcP]R\D]Z/HMR=FfVff_bJ=_dd.BZ68=eOF0V(AE>g(EF3Y^C:YMHZ7,#T
94f_:<8^>GF>#d1VH3GJFaG&992<c.GYAL4d/fY#V^V_+0LS0+B>bFG>VY5LI)fQ
>eV0TJ]GHSJAO_:PP/.g@73eN.MZV0Jb173N=fZ@J#(3Z1fBeA)):?)9f^]>O[0S
D<0)JCKUUFRF\TG88(XUJ=,0,7BZLMc^g+-KJd#H&5SS@bI>C6g_A&>@GO5O5V(&
2<gC1@/6Da:,@eHGdg9#TZ_4KOBQdT=Seg3gH>8D(787];0g+R<-5K+736\Q8[a+
,V[eQcaXVXLUdLC?(d1/G.&YHG).0d;^.7P?XJKe07W\=,/-VSO?5)A(Zd]S?6.F
E^.aG1:U2,f@5J7ecFa0]B3WR[DF3e3V(?K@^BaAe-G:W/M:AT(GDIgbN;>T9R4&
1D3?f,EEQ3:P1Zb[B?a,9&ROH)OI6cV3cUd&M6eaDY7RX/N4c6X.:gDg?DFO7;;b
-a4_LGDFW.a:K6#97Td@GXR&F+S3YH?KZDD^IdT:@9[1H,aDCQL^A.BK+.a.f]Y]
<JOJVWgSXT3,@P<_-_@[I)UX1]5L#9A@Y>3XY.FDeX/+W\(#-3RPeJU8,-UHKO6d
CPeKE;I#,G7(YQGY?;<T,P>_fE9-.DM-82-+V@;/7)gL2DJU5?4:X<SJfJM]E]85
8>[3g&(YcTMGY(K2Q+38gQPYTYY?4#?X0c#1)[af;5KX.3G^fX&G^P.ecgd+V,BM
2cFC8CN1/8NZBI@3H2D^c]_H_GF9Z(IQC73JEVQ_V&0,VK8&(\Gge\P<UG/AEY-L
Q6:#Y??M7,)[KYPQQ6\2fB(Uc;D7.G]7LfU5)A_OS@AWe+;Ud^R8]N25U(cF+gd=
9;,#?c9#Q2GL(#Q31>#IXC,BPO9?(0HK=2(W7>Y<(<=Id)WU8;_KLd71)_bD>]95
^<McPKS_+db08<M,EC@\b9_55cfPZ[Hb6H-fFD<UY:(1PXQDBU&QaPF^#YQJ^3(&
5C+;TQ1#5V>:&Q5E<&B,<fREQ:B#.Rc/eaI9e-@T7O=X1W9[?J4[\g3IfSZdF/0R
MdSLL:.J-fcGBJ<@SNBB\5HGZ^e2_bG8egA:NB/)Pa.DM:a(YX,.;^g^-(V(?6+/
O5\Q8JW-I.d8@M,1B)A_R4=:@(_>2PJ=D<45DTA8Q3&5=,>JNa/JM]TDBde0AVAg
>,B@,X<<\#6IZKeFY+4&U-1,=I][PJG,/>G1.T0KMH1a+5bTA^3>=ZLR(4<ROOPc
-?CV:U;O[W<d+8(E82M:[^)MCKYA#-e9<8b@JR9>/2WXeQgEIN=f,eB=O#aPXH8G
K@M^I,8P^P>OXAKBV,N[7:3a4[#?CL#\fcU<E2V_]G4;Dc]UNZ_[#/)YHgR/WC+Y
Ec_;F[YM-KN/)G]_>8FWP:<.>MKd#;2)&8),]CQTaNC]8U0L-Z@7^/2L8QDAERBM
?^4.YQ^.SNR9>fQfP8ZA,a-P\;RDSB#FO8ffZ(c9AWH:G^TLcX3(SOI<-\1E,2;U
MDXYTNG1\bbd;,0<NUaH)_UCH-8TIDEf.7([KCL>0MCbc3BX(6(+/<<6]\HB.;=3
Fg_;=B,7SK=7G8Q<:.aG8715&S7W<-;?+@4I>f#FLJAYZ15V]<Z^D5X2N/2:6FKC
1.(MI)90e8B@K47BLOL\,^0>0<@6Nb[\#F[@XNdfTdTH.N9eG270),):3MF=0BD[
1;F)WB8NE:=\;XMA5_(_&,Ac<@e#WbDUVQI-aE##]PK\;?)-,OTf@Y:60e,b#-g6
9OZ,<0GPaeETc@Y;HQJ678@&5?IL@=9b>B\7/485If_ST.d1-bJ0Ke/-D@&6X_Y5
;Fc.D2_(R^a/6FM-?2gf7.ebXObTdF<5M=PaC696E[QKT9fG1A\#_,Sa^>E;S1L;
VA[WJ4dU>6EP3b_ge;;g^0#W3\6X,P#Y7\aA[[K2=cJ;3Ad;GH^;=/3O-IeC@I9?
bC92&5QJU4dN)DOQ6WVN(@V]aN/U>SQb\TDaAE@eeaD/VD@F=TT>2A--ZdGVQ)R&
)R2G:3AN?9:M^a2S<W(F9P7ef#bO=aadJZIYR6.geS<&HY2d[M[]4#>)bgSbW+gF
&^Ie0HbPX+JQ@a.bg]7\A,X5W2PI:I-=FI_;N^7gSJ\K9\3_AP.,K.HfW?I(;e4\
/L:1,<NVce6POf>,d\>#e><XM>A@RC16+/]f5]@DF1d(8IC49&5^Q@N]70Z?CS3N
&;9\GH:Wd9C65C?)J]+R8IH9Ea]SE>gMf1WH,2dHCf:dGDJ+31Ya+OdgP<8ZgZCb
7B4A:PE32/OBHL?KJ+4L2&^[ISR9M(-_D2(SUFTGWc.TXfJOCfDB:G(I8JRSF@8A
H1A1O(6P91,\W65=,1K[JI]Sa6E>4N/3UCac=NI[8Y6FX&PC)3a\\OI0MK@GO#&Y
;f=7:+@A+#EPe5.<F>[.UKQddL]X#MRf1G3=BG=O2?U,^BOgA5LH(DONR6>J?[e\
7+K3eYGKLVD228W:X^TP1C\;?-9=I9Y:\c(e85UbEI]9YZ,#?1S1R.bA>@2/)gMc
eX1D_gNeIJ(d)A]VWIH0R+00E]]>P=,<=Eb8),NOLBKX3=.E#W6ZP+eWfE\BTLJS
2)X>Zf26(TSXDg51PBIe?8UHUCKU.]Nc?=]J+g((9]&\2(91+?2=^]P/C6aPAV>I
.7,Q9A&]/1cLOM+-[Nd:g9SY-;[+X6Pd@-VRZ\G_eP@\dbT>1UWgWN2<I>8(T8TO
\4bW7/8RLG_c(eaLCZ8aZYf;>J&@eZ+K;:6H(=TePDeG7N8a77Q/&PB0(P(g@F7N
/R7#1,c,;^)cY)U4&<_CJ<Q/A/+<Aa:DTUEVX#0E^ZG6g.YJK;3U4#6^NZS29R^4
@G,Sa4cXDAT<@>CBdM2CI0>=/HWT:T=DRV7DM6_C:>F(E^D^R6SF2IKT#[QAR_]-
;:E0PJ^Xb]B>LS7)X;8V8S9X4S0a=VXX[cE<D8ROO.=JC3=BJ<gCKeORCPANX-)L
[90J&c98;-F.X+HKU\\Z9)FeR(#ZHaEC\7B@#B2CR,GD1-)BXYT6gAJ4IB(5JfN]
4c_c1F]M;:F(AIMM16W#cV>U=:V86(+F@9R?cXFb9(1OS6&91GE0#D=Y?M.F>XPW
M>RC+0VVERe1\:C5,/S6^.ZeH<T/3-g[CRdD0CZKE-.:;5,]H_=\7T<1dOfB/AgZ
[Pf:F<f.cfdL9LP1&,dS3KdBfc#Sd6bJ<b6<?eT/CB^NE2MPcY^61fFR(a6GB5XU
3?GBIgWMI.VR,7M>;J:DaC/BDZ5Zf_ad5d/@G<?4N=df\Y@JIJYKPgR6P:DC/Q;E
G[/c1ON7\KbZ9(L&H^W2T[-4O#J?61+>4@3EYU6LLQ6ag4D>_@:Dd&OQ>e6AfLfG
R^,eS6F3?&)?&5c=^e5H/AC+D9/]/g@+,=3P=2\ITCO_,>9SH7ZH/c&VCM@OFGDI
9G:U?f#U=.\QU<\B7\a9&:AEU9E1(V.T9BFO;UL1/:B9O;fN@dXc>/3QT#FT:Y\X
SORT0g+Z6Mf_C-OU3@.fT7fdE&)42J]gE=.39-^I43\0:;H7B0EVLRU9=#GAP6:;
QG@4Q^A-<f9CB+N,WW&4g\O+?W@4K@N[BP2?.GTd[HLRgcF3cWI8ZTXgH_+JAGPd
Cc5F_FIcaX_ENCS&U/>Uf;XF(D.<GQIJHd#4aHZINC@I[G\edMQMPTFS:EE@KHG.
VAcY-A2<;CNUX1#M;,Z6NQ]5U1Y0GHEX=(_4ZVV<?bO1DHJ_3gUSP>J]9LRG=f63
\fd-<#a6U1.D621_(B\(g&7_/S[c\E=D:?g&g)PB8f6W=b_T/8Tb:9F,0[,DLKSH
K2^_9_O61P=g[T-aZZW?W2EEf4SUL-SaEM/?MKA7\fU-[WB_Q1ER;-XKfSS+DX\:
_g.5-/:OUa:6_P&QUg]HRa\YI7K(2TI<5.,NSSX^)LB5c>FX:R>L(6KQ&OLS#)U,
<LX-#2#TXgVQ;0ef<=0>INA]_+?0=R@A>78KF68Ie[#ge>(?Me[W&I02d^(A6CYP
-<LggXC)g7&1gW4#NM<F,.@0_W&GGX@GfFZZd5_[FH.Z7T>\))D:(7ATcAaK-RYN
PQO0UOCC,>OOa=U(WIgDSZ)L6KB<5DI9>I6e2X\B)WTN7De4;(EBgDVYFL,)<cAe
+3Y#<)40ge.-U>:[a45a(GYH<SOW2e9QLbfRXH556O7#4ZbM7EaHTZ@,+S]-=\L_
@HF4DCPJW>N;Pb+-,Fb67@UDZV^L\]TgNg8d0>ITZb(MJ0cZ7RF:(dW?UZ.Gf@(3
BeCgSL5M)D^FDBXTM/T7Y+Z3f0\9[+f^cR[g?2+5)Y:<g5IM(08(7PLUbK\]FHWV
_a?J)2?<Oe]F9,U++@=+L.@OC)e>[aRg3UO7g]VX<XF9W(TUB3<>5:Re2b?EHOcC
K#;L/M>U,O@fb76F)fRC6@<68;Q:a1IL/5#edf:E3fLf6?4:\#bcF,M<TYe^<g^R
a--&S=BMVeN,d_@=_)/a_fI,SR4=E<\@+4Wd\.DNPQNbTAQ5G=](^]W?3;,fBX2K
C@+K4U+b+4a.XeeQK>NWb]b7:>L7+7DV0&3]fUc(0^FNbR(6+Zf[G?]9OSGTK)1(
aHFE)8dY\[Pb)CDE?9N7#OAW>&DSD]<]:(?_,.1+BE9;BPKRBfg;Xa<.[]3b>2be
VWNaZJ;RIAWb(cY2C6>4;<_448D)gNd15O\[#GOB@^d^J\71<0H#[6P\5@c]M2Bc
S;EY0>).5H2ggPCZA6d])Q4gH+81Xc,J#:08Fa1AM83_H)0KS[NHP;GY]6?7K\;T
e7E<gW@,e_J8]SJ3_UeR8QB<WMGg#@=^W^:@UY7VHQFP#0:\BgI^X(K&TKEWS3_9
<X>QLU4FJB;KO_]3WV[4Y\/OJ@a,c>UG)P0N:>FBZD;S<FdgG+6YX[gc)fNd#7U&
;6dV-=O;QH5ZE3dO1aUW8DcU_9<<MH52E3-JeHbZcT^^W1\BX?+<551I;8\D-M9G
EF+P3RY,OPN=&]0MU=NMgR[G#G7#:H:2EGO\NSGB.6:gJ\WI;(((+,QW4RR)@(:4
0S)f@gD+5>e^FcfJ4P4cYaH-E<cS<,@^.]^TPOEOU&:RM0B+>ZFQ_^A]7BE<UJYd
@_WOMX\d;<_G3U#[<WUU7bU2X4K,F0[0VfF2ST0?&KUSUa.[_J/B?++.4A):.JIX
2FBWS_(&5LR-I&PS7_JKR5e.IJ7cRc&J;+\A)cgXWO)c:?/P<<[]e<[:8UOBG/T4
YbLdJ>6EcX66J2.#.X5abUG43=bOI=V2eR9(=H)[Fbe.(XgFS2E[;g=XbR?Z7C7_
Gd[U_:GACU&H4[#W7YK;/c2Q(gPeSP&VW+LdVNe<])B3.5O6f:YFRPW;LcFWMEMU
3[C,>^:6E1IT2>,Dg88?#b3TBOC+TO-B(gNDYSR8H\MG[cV:-6HU^S]Oa9C[W.PI
A0H88FL3<N8[V=:df,gQ(K<dVPg@Ka5F7SKKd0(a<6d2#&PFK#H\<4&(\M[WHc5U
G7]3)geL\L)=O[fN5\;:FEZ/RU]VVAQZXaV4,F:O,#7#5XQW8@VdC7Z11/3;d]EK
^I_=F2R7)dR7G&f_NJ6TSeES<T];&+9ZC?ETfP[9TPP7DeR(UeT@Z_Y/.HH753,C
ZgEPO:E:.34;E.?XQHNJQR&QA8W]2;PfG8gX-ORIN2>6(EOHY2VM@[Cd\3<@L.(;
Q::-b/<g#+c]\WQ+>@g&>5J_J^c+gHF)DJ?7ag>gabI,gaP0VeI1=8SZ8KTPeYU/
eA2SA9EEfCSP<W,;HXUZB?9SQ-(]C/(J?K&Wc07)HE;eP\I2\WH^)e>#+9P:VTfM
7-^6eU>KP-#SHL=1-JHJ_+\I;?O?Za68(M)PTZQ-UQ7a.a^Q&Z;dVMA-7c-3\##a
;.Dd=2&V9a<PL,d;Y=c)WI>FV_2XYJ7ZJ</bg0[c.]HEb&H/K?5):6O#>L[SWCdD
B0D#D7X,0b#0[c8e]c(YVaGfWgDD&SXRN9;TP610U@0\CG#X1NP8g<JL7<&;^Ga9
Q#@R65DI0=b4;fX#K@S-aME.1;LD0BK+)+c3Cc2RIT0dMAc/X)I9=02M9U8N,IVb
2\9Tf1SG:?.AXG/JXA9?LD#:?FO/M8N^D()P2ca0+^+62(Xb>[?WKed[f>:d:E#\
HK,Pe_LO;08dWJc&C@YPY<_;:=dI-5d3B5@&^CO1eJ7dHSA8W#47G1OZ4SaW]>11
@-C>_4?]Z3ZJ_@?T;X?,a90^^P_;)ccCe&A.D>7@dL2GDR9:JG]]]g5M_LB-L^@[
3;W4TJ]T<2Y4eIH7/2aVQg.LG^\=G8.G,K+NXE^5EXQBc]5LC)BNL]Sec)MD8dI?
^D>N)L5Fb55=L/W.+OV(4M7<I.;bYAdT79]Hf+bJ#@bWE&>:UfQ305-^6Ke+,HJ6
c1L3gBc-S?&TC_d<I9W(1H(.+L8g/G;Dd\A8#G&2;,UfK/U#B\d[8bYHb]f73E5Y
E6NV?QQUZR5e@@5C2aXF>/L<AVSY;OS@g&5@3g\a_g\H0@TKL8@+fR#;UYTbU#,(
J684JdU6YHFDOc9/[g&XbE&X\g1?NM&U@J?2RL0=G:Qg7?4:9()=eW+g+.-W2Z[^
1R\O.@.FcY[)6V+P,]9.&BDIOS<;MQ_7bPc=^K?HKKL3Q#[K;&)4+U^#VU3S.Rc]
GVf:(N)ZZA4PY^a4YU=W?6PZ@\:df8eG/FX61Ce=+_E_A;K_WI&CRSB#Y;4VeF\^
P74BJMeCDB>f/[9Cd;A<Qa>>[T6,MAGNeSNX&<H2YE7N8-_1fg868YF+^5>DbP+I
fWGM+D[g55P2&<+AT34J6-U0X4V[H?aE?;P+K23ge_:FLNTY;&ERC+PX:PM83#^/
]V6WSL)Z,)OH0#BbZA:L+<IN7?U7<QFe74E_(,+ISL6Cb3?(;])L_X#<?g]@AE+9
=72MAC\P2=[T>6T[;c>U?d^R7b,ac;FAdVC?H<1,^/a?[VPF]N:dM@SSb9IWB7B,
g&_<ZT/IP?5Q2]7M2dH-]H4b&MZbQ5I_X./d<M(PI).XJJ(L1G]I:6.&HR;@gDTI
JR4g9-W_R#S;S=#/<b>.WF\KUgGaHXWPBdZ8(MSa>T4W0L>+5g&b:^A;dH##aYdD
&>-DW\_^U70TD?UWgID^b7VbA,ae7a+GXS4O5SA\X+UZSdM3_R5e)SJDR(>?LMD5
dKB597SE)(+,a8@g#OJ7WQ3+_7PKO3L+V,-(fF)g4,?GSg/c=\WbF:JaUH817\Y-
e)_/^>&@[W[)bHRVF?I6eF7=BB6\Q-HR/-F<TVI)1;a]8-9][P>.HTe16]c/@/.D
+0,MV=Q(bR2ECYN7N.B(ATBc)VKX_&d)<5C=D&d]1cXCE?>H;P]6O@Z?+FIQG[V3
E]:D=9V-Q8MOfV,_Q4FL+,-3W[SC,9OA+@WYf6T\]R7XZ)?4N^-+g[)2>-[PFFHD
QL7e+7FdY==BM2/LC+;Pe/BW95SX^5Q&Q,ABXZC/]A?_J(FZH>WUa083BQGW-(BX
V<Q)[gD(A_CVf1-GT_d[DR>LG+J/V1KeXVS7<7D1d>G0;4Y0e0Y4e.UGGILHDBR)
[3VRH7#V?S-SggD.[HJc1H]QJ6;V:g3BF70>g313>FbOS(=c,eJIHZ(^:/Xe;RSC
7FQ8]A-^.0=&._M?64.08=Q,c\TId)a@I2@FXY/#f1;M^MSF&(59+/[EM04@.70c
\9GUL+:Q6&,C__Y2(N9R&GPE2Y6bG[BMa#(GI,SS@,D.THd<DQ>RBF.C&G1.I#9F
13@B2Nae4JI--8?AE?C6e9I&/SQW@dN=HP+@KcVYOaP;L,&dDeBO#_)43a?b]D7C
/gUfXdUEf2A_7:[>0J/caECF#XeT4L=\DCSdZ2cR\Y>/+:MLL<SS]=6NJ^HUf#0I
cLFMY8gBfO098@@AfI.;2K#XgaKdY4eR1,S#,WK+cN[#?,F^K-P2J;_KgYX\NZE/
8XBPL7A,ae-87N:H;^BN]&d27P+V#b1Fe9]LFGdc;Q^a=++f;J0bfD&_eFXV::P4
TY16MM6\AZd_8@;JBae:7b?L2NQ3)9]M#fa)f)GQb43P=b-WEBW>J2Re?H0Rf1ZE
SC\eD7A@UN]5[8IK[ZAIOP:=,O1b1g6GEKeX7Xc.bA)DO9^ZN/Yg#^TPL?HgL0U6
a/T&[K7d9E[Q85DX)H^=<(\c(Y=RQ;QO5BA.06\D4aGSP9eC>^ZRII)JT)?&GHH9
^4TeJB\MI?C,X/3AG:R2D42)8GPU]TfEI<DK;\)W((3VII?O7Y_-OCeVI6Z[\>]-
gL0fX/d>4K]+Cgb9\fb7[W^Q&GN0ATS:9BV@SQ<UF#da31[7KYIaWa;)aES(CJZ<
Va->75N5<1#54=E99(U.+N[>@V-4H]7ZK]S_5W];QA;1G\)/0^d1EaW=^L)=CD+T
9bA/FdgW&64JCS(;:1[V<(Ra59:>-M/KRCZc)<L.MH(cGdG.#>90(+\KTS[/gQ)M
-[P5KaBLC-Y7N7OEC(e,T\H5;b;S_H8bFBW5BIXBYO^P9Z?GJ912\R=80AG7=TZ>
@0?RHe)aV:4S1e)?UNM?cd]YSRFP8,a&Pe)AZg>+O/g]We^;(V>4YI&X/U_UW4Qd
5S48^15BU0dSI(9]+7bD:?A^#Q#01U=-J9[P?Y#8L-QULDF1M+\a:0S@RYYcF3C^
HR;Q-LA.HJ+X7QOR#6F>XfOCDcBQ^MS\OWT](/@K,B&e?@JH8gBWEQKf67B:VYe^
MN+RYL>\?-PI@=O^1CYE1:I9JU1cC69b.g0\?87ec([WEe80#/b9R(NL<,/@TOTA
8;<KFK9PJ39R8KNX[/AWWPc?QbHC_,e=&QIe9CB.@JH9B2G@;#:KL<[/@0L>S>08
+\(F\KMdITA[25OLO,g7IT1L&<]1f,\<QU+UF&VF6Af(0(PbQgU-=>E3-Z5/JCAc
@+-7aN62_LeGc<X&D\1P;_3.M)Q&Q+XaJ;^<]?9+4<EYbLMWJgaJC:cU-A#NeG@=
Xf=g#&@d2/a1+?ZR/HUUI)H-4PQB&QdD=RB,E?,F07=G=+B;GUB[_\B,?9b,aH8V
<OKJ?041T.ILEc7YE&E_A4#F#bM:eH.6^U>YebT756DJSK650cA4CJ6?-K\X)A>d
S4)I&A05A0Q&A.c4_WTeS^2@WJb>1H:QTU<eSS4Ua#K;BGa&S^X3GNX(8S>,@_4:
]@117<E^>b+3DX#ecGG<fJ[@D7(^+dZe8F?C\BOM.aUc[0ELCJd?aOL=N<YL9g1W
]Z.VafcAFRO+RHF4_Q1+A.B>1-XbG2)gQF1a@WK@g;RbTCRJ/@K^4GGdTMJe@G&P
>b+NWQK=A_LUGGCWB9C\C:[<;3+8_QKJ+^IJLO>62BI^D,D^T0R=fUaE&JIZ,2g]
gH\eBSUYa:_#S-U0Z^[;LaLZI\GT^&K.0O?V&]6\QF/+Q;ZBceBW[/X&#?2+2K6e
)GD.BT9BdC#DG,EX>Q,T=//6Z(NUT+0Z5(Z-EbC<bTM74<CJ7c]3L:[a]-KCae.Z
WI<b4F7,gZMZf]8[6=GYCS>OKfa+>#^,AS.TGW7VJBX14O#@PO6ZgA(MU>c,UT_6
=2e2R\ASTQU(A8Bc=dW==#)Ag:7KE+V6ZN&T;IE(RMB#-eF<@<IY<J(A.,KP5)I:
e,[+S2\,@Ie;:^LTJGe&c8]:3Fe7OfK.D+[I])3=8#C_)D(N;2HM9&P_CZVRZYT<
F]]Z1fPCS<&H>-2WO96][Zb8.c(]=]T+O>9MU\O,=(K4BL;V1Y4YD6EQ\#0_AWO@
;CKX2^:AGgTefcU-#e@\dK,T1^.,UOL:1IBJ]O,CI_HaA#.UJUD1JCYZ7;]&Zb/I
<gK9?d6>MV/;8+4(8PgML.U6M.\cT7L^6:,9-bRNRa1QO<NY[VPL<D7W4T0I<b<K
P\c@d\.^?U6T7E6G8M9&Yd0,B+U.-.&WMZ@X##K8B<<J?Mb&g32A8P^@e<N)XI3S
QM3g.8@KH>1&;c]OU-YfUfS^6DGN8=g-TID5]/cY.OLcTOX&\7BcP^EgNf\4@8I?
CDO;4#:\>ab.LAE#RSMLP+420C&]b(a^_XDfCI]PT&61<e?Y@+Z+<KST;)f[cJ85
+0^N=30EFK.bHE&.N,HUa/@<H7He[3:1a85;2/?Pb-X2fa7MfOZa#TXSg&]P3(1^
Q8#@?^].RJP;OJ?Kg9@I+cJX5SF9WREM9A>(YYNc>df--IXb0Y1)3GS1\RVU^C(g
(G]1P,G^TN=TW/[OQ70;&^e:S/5H)3E<[GBfWcU;O(J#HfF;VC+]Q]V=5TJF?QFX
-Vad1gM,.YI?-?53bX<?2>_A>2G?E[1@<P3e]e-<0VOdaRSQ+/EK..64;fY,b19^
DN2Ua3DDd0:0/P6M4S@DL^KQ=TE^13<3Z56cAP)94#K(Z3AM95T,T2YL(8ef)\+7
_gQR15H]T1Q&+N6X5:]8.-&=>g>@d7eXLQYAKbdc^fW/EDS>e-,84V\gJA;-SBYK
IIf.Y?cK6^e121f32)ecV>IH^W8CCAGZMVD=+:I@I@+=\XH.+2M_Vd10@g#1+IRJ
I=LX7G\X8ODFa\RY5A^OQ4_/fae3AUZ87-TbFM,RHQ^(>S^gd4a1T_Q3:XK@>d#\
VaPJ&e6Y2D[3ZS3.Gcg2F.9MW\>eE/KF\U(;d2,[G^I^TQ3&EX85beNYP+260]X]
dU^Mc8<Q6K/:GfB>A;2V1e?-P084eYV[67_b0f+&6XU<D\RF;a7b;P?WQ815GbPA
9?cga+I?WUTI[YY@PLE1V[Jae#OJ_R:gQCR_BV4K^FAELQ0>b#^USI,9N/YC9_?:
9e8X_:4&4J4eB]_9):9gVgI]FDdKMT6LE)@KX?QOFY-S6]G<&++@F<ZJE.[PQ5O-
Z]1I.H/:Z,f?C_<-DQ.^.:IS<3fc[\\++I)EK5O/G<:Q/J4-KLFb:FHg;9?X<S)L
=6ADL-IdA[6D4_Gd6^9F24>)MB>/ZHO6/UVaf1b^CIO(4E6LEOCV-(65c,=Cb0F.
O#g6ZKCXB<5G6[MY@U&-/CHR5afTfGfRfWFL79T_@/TGL?8W[SJ\,@<Q.=PQ^L<R
;d((P6-VU]6NNc-g@>I<E;14Y70AaL<7:N_GDXW_QOU1&.=R35fd#JCHBDPO+aa8
,6A6a_^XW9SQ.XaG]V@MI:)ONJVc^MRYEMd)CI(-=[DfLBSdX:^=fVE7(e<ANMK4
E(TR6SHKYWLea<7?)8?)XKJA3(,R@VLT=H=XGBg)_#aP^#W:]d]gZZ[EK6ZC&:W>
.,OOA0XA8UKDW]Zg.3eJU\S[([a<3)d:M+Cg+8^N)+NMSK+GW-DB&aSN80@:]Z]^
MNQ@VE;T=9V,\8I(1^TfXC95&63(.:U<P@aCO-@:O+4<B@SSG)/+I;g1[3SZPMRa
9R:,cNVBBf^Z<8H)e7_)P\Y^=[UO8GQ_JHEM_S83e-bTgSWg(=,VAP5CG42c/+e3
MLXXATYS=6LH7)DTYZN0bAM@T>##d^^RHLJPXG11Mc6d#a)7O2V\A)WGg[\VID(_
S<;^86_2&;JWc;W,R2RS-&+G;PGd)gMd^#DE=]O;6-1]#CZH];IHRK&H]a7f^YA1
YQfeZX^CY)]_[JDL?6JeT[Y<56+0;L>2V530Y/>cERB0GYcS2c6gE<2YQg_Xg7X?
dX;bXZ=K/gTc]L4E=\FTBT/I0/PZ^?ab&C--V:[A&=.#R_-^R)X()DQ=+K>10VI#
);84G<VX\TLH,7?6XLC2a+TW?a+(\-?aeW,P#Yce>C4V)d()7^T5[Oa1[eWcP33^
Q1#5YeA+ea0,2X9E.a\fHY/16f=(c_:77cIW,\Ea)2IbJ\T_XHY(GIMKIO8OD:.2
;3ZN1/:0CgWRD;O\.K6eQ4Id7,5,#d@U3Y,&\Y8DVG5<N.b),:>352R\<7J:=O=O
)V]@^1ffM6M)c[(@A@f<<C_[c6B7.BF=V>,OM0XPcD1DIa,-/<dB#D^E&[4QR]J[
1Fdg(0^,+FXX?g,b):(VBZYTZd5AC@EJT1-&dW^USA5O^:BfVePVJNR&UV/K57O=
Y9/GZ.N1TN6FM[S_6=5L.32PL[gD@N_=HRI.<6&R\R:Ud/FO<(PQDA#MKKDRUc>d
=;T>Sc_Y^XTL4bHTDLHOGc.-)a<-g.cEd_-gM:31:f\RAO>C.f[\.?ec_N5;759W
Aa/M0bR7OTJ,:S:Ye2@_7GdDgCfV[)?;Y9RN1PXN,4N^Je#B8E&_Ef5-7_O+g[6F
&#Y([.;R=ZTgNM6/ZU\Ha8-a.<+[.TDOMNaT3I,??G0ZVV#5QR1RQLdCLRNR=-6T
U=K(ZH/Y^Dgf3\WE/RS]c\0.D6>c=ad<@1+X#f0YCc[<^[]V?Mg6))N@;Wd^VO;T
\;KT)@.I)FP=BLS@3VU4Ca9=J2eIg7L>OZfDc]c+92<<Xf@&LS>\[\>Y-SbfN:_Y
M;<B/:N8KO:HfK)9.-GTXH^([LDfD[90gSTE8<5.&VKX8Z\74eJD<[#a?2+@Z:R\
85TH:R6bTS56gU&Sb3C.HT&8SC&9GS/?AW6:;K(YZ+E6;ccG\NW;^?\Pg?+6VJ:[
D@U1aM(0C#HQ-U@YA>G?PP(+c4KIKf+PF6_RW?XL^6VYdL9>@E;RO>E.D.OA.I5I
O\/RfZKZd.KWL^f<WG,2^#c]/9J_g1\G26:GIe5C25aDT:+1e[6fc8>5.7eOb4B8
)Gf==Q1\GaR;F.QQCI\E6Z<5ZNKB#SU[60M_BeJcM]\Rg?UU-C5b0(Q>bf6Uc.=U
e]d=MEbQ(C^2FW65:JRC]7MeG4F+S\1.b-,#Wa0(8a3://]H8M>44FXBD)g;OF+F
4cEe9FaBIggg8<)^bA7IAWHJXVV^0=&d#\>TG3#&,YdgC)/D=^]?&I>8-?K+\>E;
MLF^bO&7#=789b)AgQT3\SK)OMVOMG5=M0<b\XaTY7Q4.V[0eZEbb9a+9]P\S]a:
d7c;>K/SA=\(>1MH542WeG=,N8INKC5REME(acD9O13YZ3WaC.C7(-=G?DA36fG?
g?3V1Q4X;V2[CMKBAJa)Ma&F>28cWR::a##+H>#&\@g-,DZVP8H:#43S^Xf#POd(
FbVBB(e/9)cKUI&dDb(Pg9H/G>?>5.=^LJ<9R,)RDeWYE1c?PQZD-/Og\/gF7WbF
<JbOQXf#f7=XAVAM<12]5L7ZZc,NI>\7A2ZIG>1OCJ=WT/-Pb5MLK1b?-bJY>N(J
3H)XCK.ZR7gVX9MA_:P]1DG<AI;D<cDVg@0&C>]NY&5_#,9A36V<D3+SaUdR<K#[
eVAObS?X2:BFLbPf=9f)\)75UIES3.[\(+D/&8F/1IO@WI\ed63+2<#Ta@<g._^F
[\Zd/R5BUZ[;V4#:<&I:?]N>2A5GDKMCF<Q)#3BgA_11>;^Q1;FQ]I).R8E?A)^5
Z;CH7SC.+3C4VEg.3>0cF?P,WXK_?0K:Y,W&#K?FX9]Z]LRQ?caI-cPFQJBbEaCM
ASLZSAR_JWcbUH-IeU\>G+dR+[6EE=?\41JADA0Tg6>F5eeN<2\RI>,LPYfE<944
T.VO4IW3?^XSD-9.GD;:Ofc=5\Q<a6:-e)C]\b2SI?W8#Ia4+6QP0@?+Wc^<WI2N
a3(SM1Z^FXCV1RJ?@S>/R/8(b-^e+&A6<Q#K5,bbEgW\UR0QJ[]49U&W+^bG[#,=
3S8XLPaD<ebT:U-KT\=Z;bfT4?:Fc(5TDI#C-H07-?.XdP+>Ke[FO4UFKZK6Cg^L
=\.8F?3DR-@H(NUg=HMQBdEc<R)e_-<.F>]9?X57BQRL>)VN8007AS(_]OQ+[2@+
.#C65X:NOFbGe#aKZSCde53bOP,1\M:)85XVER#7YKYb]N3O=Pdg/+;G/f<,F])b
3JP(eaP\;c9cY7\XC4Gc&=[f.dfAEY?):K4O=A,&/b8SA0K6D?Hg9V21g\EJcZe\
FRV-E97.&R8#R1K=.@P;FUCcT625OJ;\(:[#_3;Z76Jc08<&4B8NDO;^32c(DC>0
C0\(fVgJ0JSd2M;5f>+/aFQIT9P19QF&Jc7D&?g)#_.3U97THfWF2VQ\<0gO\T-A
,PKB_(>^)=W:QA&8]^&b@g8+.WPc5G0::8S9#W+T3Q8_e;5:/S1GX\I<c-Y-<7a(
?J]AgQ&9K24[QPaN#SR?@b\VIO\e//?75173<,eUVcOA3=;D@C5f,3-0_;J:2B(F
2LZ>;#:VS1Q;\0C;g-L<JKC8Z8GXWBece60a_;#Da^J0CYFT<E62I-8b>A.RE_3<
P>M/c;,BeM&:KG4:5)UK-EIFc_^1X1XE,Ba\DE5M;?>Y?XC[?968L3,7P\->6_)I
&<?4Bf\JW]TH_b][#XUd0I3B;:83\0+b1(R1-7>RcN<IZW)de6([V?WX?.M3OfX8
/LMfNEEZfI2:YV,Z2TLRV/XP+@/ZT?-O?[&>\P.U(M^(?&U4CBQU?YbaX94ZP0=D
d25PGD8IfEd4S]N9;_=eD>>:29DbHK[4WQP._I587?X0Lc:Z;a?O1JE.EfYNX;ZU
H#/Rg-DN1X?GM]P>?WG6YYd\QLfMJQCIRP^N&[XE-M=^QXBOS7+(7)^B<Z+M&c[d
;7L:4WY6cb.(c/;-ZgN6,5bT3G#,FO_H=L+P.>Z(@V>aTe60Dgb7UVBXS;N4aE^/
38^1M@Q:H/F8)+WLQ\F.&0H@H/WDHI/aU8DBZM:M<J9<A89HMTW(ceU#7?g?@aY4
Md#:O?UV(@UQLHC6P>Ib5ARN-GNWQOMGUU;L49ND^.aN9[;d0UaY[2aZ(d\+G2eS
OW\V,1&B#ZGX<-KQ9IF;?DLLXJ\W0@Z7E4\5V:6YI429FCP\&IGSL&f<=<24.44d
a23g5(E@?GQb+Q;3b[[fMd,\F+&.LWCN,cKd(G\SSTT<04];_&<^GUYV0S8SLT:W
4Wg<6AacKcST#VP<[_&eV?8b,RE8)[V72).?5?5C(-L16/QbeTJ2J6E07DL;@JF,
?aA:F+3YYaa1.EGaa8AZ,JJ328Y/)c8=AI@3Y0>P4^c[>@.AAbS8F?e@MDNOS[^C
+bZ0CF\WF(cEWC3SKL(JF#PLd6<08?DDJ@3Q0a_N2WaS#fG.LYPECcN?IRYV+1B2
/5Gc_&H)-X88N88f(>+6g<^f@X:K5WI\12<2[<1<,>&VJ6N@:9V_[Z,:9E)O\?81
E[FFWe(NE.eFPI:H:gT@CYDH[@RUb?)GNWC?1<W/a\PM[<,EYc+#gI6]/8PNEHg.
@5H[YBR2I=f^HX0>RR,JG@0XD,P7ET:/E]<X7SOa:9TY[fGG:bGH+<]GT&NID(=e
aNdDX_4aNI?fSZU&L#>b8R:O-fXA/+]B:6MTV_<M0I413eIM\a0^LeYWcH-K7Qa@
7OV[/R4@IWD]7D@S33aW+ML=.VV);IK[[+(WQ_Pc@:G2&Ie,b#6TR.)<?=1gV61@
VUY?<+JY[7d[?_GBX.@FeM,3PQ1e8</Z/5^^^ALV;aN/CI2QJRIeWEI)WJ4X4f\U
_FU5:>)0+70YJW<Je@bXRDGc/EgH+XTWf>NR;Ld7-TW^g0dga/?UDUQHK10_;/8,
+9/a2KScK\QEL\(QHLLRI^P3baOC@O7_)+6;gHcG(YH##0<]I3b>dbLS897W0-]M
#ZMSd[e+=H\=V^;KfBRL)O7e@55[TC))\a;@?,)K/CM7F3GBW5B4\?8GAX_PeDfF
5[b1#7Q(2N0B2+/?EESSPXU^L8gKPUS__X7.Y#Y2U?0IY0;3@N&2_H4\)g2FO2_R
<R,gD^e7>X48787dJH@+@:>QU0c](MW:8KP;=D:<5.NX7W((27V4H_7DOGaCd>)[
B^I[^WN(LGF7P3a6?[=D@\cN4/L+@)efO+?D37d6PC5=UEKOe,OHII>,)L-<QV)/
#8=gJ&QW^HJT>FQaAQ2DI^PYVO\WD^4SRT^Y?],f>:c7?R7YRX5dH3)V^5Z9-e:&
CG-O&,dd(IB,]WZMBAd^Ef(R>P8bO,C-3T9.?5FgUQ?.eC2FL(&2UG&22YQ^0)3]
Q1I#=D9<QQUA6dU8[_D30UJ4,C6(D3=G[_F]J6SNW<G-#1<:FS22K#LUL(J9YWO_
;2A<]4HM1RaUZ7Ddb&+ba#PgOAd=S1>Q>#TX,47HX,1UO@c[AY(@VR:/1+5ZIA.A
dWdPU8;\JSCX&G\GIE0WW),4XfeP(D&E)b0D9U.@YOFX9(;Y/3LYY[>V/=?T<)c(
F7WU,ZR9?dB=.;_@gH3FLWg&9+1,gEEN0CE,MVc,KD;1-FgYcPK0-].4cY_dP@:I
-c&(7_A)WgEHC<77+H&/DS=?dgC]Ee70.M5T(bLg)OA#)Q7S<,B_8>,Y1\_D4a6L
XB9<O[^6<TF^,f4)+Y65]UGD_bR7C;N?BWX7&eMaQ]@Z1JBIMbdA1:9P)X638C.5
Pbg^<LH-X#16V:W8?OR^L-FASSgMPdT#N/gO6fAK1?beP>8_2])R((Y;Z_<_IdQ2
d58c\J5Y>[0N0geI=c6#c,K7VaZW9fO+/YX092RQ&<_W_=K(@WWU72NIf#ALSIf\
QW-B7a\<@2DAHJf.>(]dN.Q^bN_UZKNPYI7J7.4Q8Ve]=LEL8Y#JEb9(0;[FZ_[Y
Qae-c:;+UI7,BNLVAAZ0MGe5(3;4NTZSS^DWY=.HdK/aMO><1Y/]?]7OHa@F2WGP
7\J9^f0\XZ]:-CSE#[3EX45K?0JXg+D;<&HfAO_E86Q;1SB0#Q>D_?FEgPG_3&]4
.UZ7Ua4Z-Ab]b96&GAT79f&B>];S[:#H)I:;2/^a3XGQDII(gOV(IFg09)E[YJUG
aHBSfU7-[+S:ZbK^3Y7OQg8(1Q6ZAdF&VB9(dIJVPP10HL2E;+AK78^X04-S,cfM
3+B=b6#K^@4)7#>^Veg;d7R;Y/:d>SdKX>6SV3[9NN+-a5U74gD0FYbC+TB]KV87
<T[5dV;I&/V_CE=O;E?dTOK]?dN_U(Aa1,>,Y6<MY7M)0;aOVa2E\D2(.E-VMWH:
e^JE.G9]STGN8W<BOa>T4@5HKE_))EFf^;Mc-Bc_8:+.(J7b<3A7R:1R_.G37c)R
15K?P6XfBG_b38]IeK@P9/^^;[W^4CZ.#-H#R8Y1>?bP&K8/D:g_54@HC5UZC?]>
4Ng4H/9W<;\\/2M4D+XK).R57KU\)X:@QI<-F#BQ2Mc/JFLXA(/G1d7BJN,_>-=W
a[U.HDD<cZZSg&;Z9PbMJR##P:QQ//?4X<\7L?7;.6//LcXcIWQe:-\0bUcG(2/(
g)E&g@-@XC,aJ<XA;Ga19^I\AXHUATGIBZOIZ+^Jeb@2NS7-:@aS[_UeV_Z3RU4c
KVD&#LUK^0H?Na9X\9SId0bf8L2\CSM(PZ\dET?8\U;Ne_C&-IS=R=e04/)4_3P-
K_OP1<UHJ7</N&c?5XA.0U)Y\O8WFeH,(d+IA,EQAZ,DKQ7Y3,(CPO8.?bM5QB\A
4=Z,fZBeX1aO7aO<-e7]D1?@)I&5NcI)&@T6CKGXHATX34AbbZ<MJMFGdENJa(Ca
YX9XM^V?7^1ZA,M1fKKS@Oad-0RQB7UVa6?;N&)0:9Y7E@SdZP\S[.4FQGKf[,9)
_8+@=d>HG#F+aS#/H+K@W21Wb-T#_[4N)C,<-=eWC.3X(5V.[fbdJ1@;;J.9E>(J
BSE1^\8@a14d9MX<e?<9ITEaa6^G&&#BKIDQ,92bXdIV+d@]E&d\b)ZSHd(LYa[C
RIFE0>KW)#cgePd+#,4aNQ0Xb48_Ce=?-2YU/SL6O+9-c=<UH,C+F=J-NDU#P[^M
PM.0<Z=a_&Y.F)LK6527RMS#+3TAa4&-M0:eY\,_/DcaW+XG?NFC])g04W<47IUT
a=V_^,OHA6O]HJN(?e-XN>^BRc_Qgg)B.56YU\c41^P4-f\f7D5VYY4d1_M9F-IC
ABN4/36\d56L?[fJ,aQ/E?g-<W-Q9Ia1gH>cUcaU[Z2OFB:044B.K<C[_edXag&?
[)3/(AU-T?T0[GRI/)C\2E/-ZT&@XA\W202;+.0EF39A0RT@\-ISVf@KHW25.9(B
2ISdL3P5fF?:5TSb>1>L@Gcce;5bQ-_AdV,MI484N/4eM0MR.N1_V#]8ZTD/eG:f
++Lc909Y.b<ZUcA>42>_B;\).27\eVPVBcZ4Jdf7b1L&>>T;N5AU\bNaZ^;ga<1#
+GdEeR?ebG<6IPMP;1BIBAMGf8PVQZZL(XY)=]7gM=Va?eMMYe5LE7gXI[POE)@G
_<(1e6X0(7SX<<-BZbPd:EPa8,8=DO5MIcdCG\_CeDa3D;e8HAQa=c&Q4ZQ08::;
GZV2A9V=3=)Yf)g+[PJ8><)+XFZQIPUR6N1>967(ZJf)QgbZVD#ME;Z.)N]25IB^
Y-1@;Ke+Xf5V>:Q+YL.I3e?dQ))Y)L72-4EK_T8_T6Hc)I6YT8VQ;EBG:K)P-[cK
K19-Ge7B63)@;4QA@::_3D,aB<7(B84YD1fR:bAUCVEc1BO\:If=G6O6Hf&fZ\O2
Pg#b&d7<KF3(Ba-a.3HXI3VW91@_T?(I[IR[M#b?NG_>)RV&1G,JUd&/@;X?7,]I
T^OF.U3X7LI]/\<c3L?4WJ3K35G^L@1CPK&7OH/?@Af[J:A2_36F8?I.[IE:?#2<
#8=>c51G@T?>D\I?43J;cA6Jf<?RH2J<JDYMU6f?&L2^0KV#?G]V302S>58-.(7]
0Ig8N0,.KC=\6N3DRP_D9IHGTQ;+NR?JgQ?YPXBd\_@T;6O9>PL7Fe#@Y_DA1:WN
f9E91dfDa,W.cXgHe9@)>Sg)eXOag)D),^DCTG5.PJ&@O1TdNK1E8P@)C8D[OC\Q
###eT,fU71[@Na:B9R\YU(M_P&]]WD@G01Z&>I\S=;?L/N7R\OU<+HeK^=c-MQMJ
9T>V.c[X_]WKcg]:DVMC?<8^/?04C#-E@[06Pb+UK1Y>c=X&eA]b@2P>-H(Y]_fC
>8gF^<3;X;Sf@S@BPfQ]-C@71BWaR?I]f(3#S)SOe)A7]<+-=W6H0+;:-)G.RM]V
[O31AVb+PGOaG7XFO_J/I@W_W8849]<<NP@aacIY]1GJ(F;<8G,U^+Q&Q/#.UbC+
BN?,&6Vde>=Z4f)#YW2<e3_;?QS2A5MPEcUSb;_b^V6Ia@==b2\9aba7XIb=eYCU
J0A8+NQ\U1PPJ.FVgdTNMWY=(/4e:CID;H)c0ae&J\#8\0e^TIgZ+S1=@LTc#-IG
8WH+Pd=[DIb7JN2H56CRM7+Dd9R=<JO.9?.CQ\bN1gNB@^Q[S8_gIb-,f2)S\1-.
Md+,O@6/P)^Y6&+cM,7-2eYX6IS[d(ZUU/J^MgWUC=a(<&agVL;#B\#=+d/<aTO5
O>6?8KEfe902:@..U@&e,TFPZ<?N/+92^7gTHdSG@ARB6-QPdW=TL^IZBICb8#V=
8bU,TFN9DUW#Z:Zf43DUO[@LdX#5C#f@]8>]#gLDVVF9=MYA,M.Yd(Qb^9IH&7AZ
GU.QXK1W@D4&6B0\I7:OC4BWHBX]I]+0ad/FK[UfYBc99^E5#5NGXa>#.:?HI+O[
+]:gd22<3[(VafSZZfXeZ+@9e(#8ZUA)+>9]UbE270aZ-).7:A68)515E8/AH-W3
5WYLg((dg/Tf0A(Ya3>Ocf4A?bGO(V]CV.f^,T2KS,_#8#bH><SI2]#1BJ<[=BFP
3TN+8VQ,=R4:D?O-6eMN>cW<]2#6R^O[SP=U^L6WgTI>N(Rd9=Y12HXYYN9JH7;K
=TRaKSBX,H(;.-INc/.NU,,RZF;\dc@>1)dKIC3_:>g7L4?g.D=.2X_)9TFWPWa:
aB/>#Qb9KVX#7Q1CEeW=UdDEU\L80NZ?T3M#_(L?QPD;TaRP/6^7aHU)AeBGR38f
N@Y+C]\H>X26f2;5^V;8AL1&KM)4cb@&Jd0bU]T7eC/?FNY=7S4.@Oc=gPO4g/O.
^(bI0^0g[PaG;\5Y7_IRQdM>,)NHRBZ>C<LE+eQ+AK^SEFe-O-;E/Y9LdO;U<M4c
9@Wf#9ZC0B1VKe1(B#C2QF0X06,<K^A<SAJ,V8e>T+B#C_VfJ7Ne4M@V2#b)dMY=
==1.F@EbgJM-2V.2DVQ&W9#PM5>CV4>S>+<S<E,A+g8F[MI+4?G>4.cUd0VE772Q
abYVgQKTV/b@\MFA;ZI[Z(@)6\7=KRMg+DCV^-6\C-5U3C[.YK,_0dS8@9Z^Y2.G
gE=T?_,5[4-NMGeUP>#TWRPgLX/.U=D44R8DA4RFX;[PT[PM1J=54U5OX\Q<6TKJ
\QS7/\@+:Y-c<9H/U,OQ9OB;>NdIGXTcW)SA>F?,?Y7^93<P3[JAVB^GVKJ>Y3+g
2ZeW440#):P>g^B]&V?,XIVQ@FIZ.J;H(QF(-JJN)2XJAHL,3gUIBJg;Q5;4M:bU
O0&W(+RHZ6^/F@[>CJb)bB^gJNL1L3[4=+9+]d4f@0fQ,UeX&V2VEK?+3;eW5BRA
>ADf,cRP/7D>7;\_#0]U=A[C<(VF39<QHX_YHZa4-ZRMOfXdBFLV#+)f_G[CN+0\
L1:fBD_7]3SLIf0V7:>X<Q6H755+8:,)fgH=][SQ0QaH8TgN-^NbaR/[U?gQQH<d
g<26cd@=a:9OdZCH@;,.KF+6]bTB_9b5#+46;UMYKER?0G2PB^0a4e#f\]F9XeaK
^K<T@Xg5TTDGQ[<V2EZa[2AA8C9b+be92gX@-H8E&3?RQI2b:BEU?UX(NQdPWTO4
.X6@a4Ve8cGNZEJ\C>3WYP4:^O=b?:f;/03[?1Y/P<CG\Tf,=;-HT9O/VX5VLJH@
EV-BYTR@<39c8BO<Y7Af&>c=aR-WPRg==8-gTDM+7XJ_;0C<BHH7>1OOf1W@N]#8
+IPGa>W_M[M<)D-X9N:)bG^QDD[/M/B;_ac3KU<FOXBD>7QR(<<c/BTZH-GKSEF]
R#?cH8DHbPB?X;011?-NBQV_,SEUBef7\<NK:gLD9^e7#=B\+dXK^LE+<.#MBR&Z
/KcL?;H3Q\=g^J-fAMDSg]b9(F=VV(5B>-\[cZOOPDc>XcV\0[CF@2A=?BTP=5PK
cT8,EEI[_FX)\\2D--ZRZ+ED1#<)1aSNT1)^UMAaUgZ[KHS0IJIU&0[4aZ3bLG5-
EaW9#+Q@/325eZ[e#-e,M+)>W(Q1=,>Q#OOPL^[RU6@Ld\CXX<eH\b2<3e;0]ZdU
;\WS3PYKJcC4A2.+FfBBV^?\1Q[XO.BPf5[^))84JF>#4^GPIONHC,:;4UU]M8FO
2B@>=]O&0\;LIC@+TE36]^/OOJ8deCNX<72,2WJ5e[&&[(5K6>YKa:2@\IPb7&^T
JRg1PJ+g=[PES^ERbPQGf3>N66G0;Yg>gGPW\ZLe&>OBab?45S>G2Ze+f=[A^<N[
<_:VXZa?e,VK[bIe+_B@/4.#:g0?-VGFEE86#N1e=W6A//68MbK.2AR;aP@[7XM3
fF7W4Hc[NK:P_V41HOd[\A&,e0-I_X29&)YT29,PgBU7Y5QC4)CGDVQN87-fV;@P
[S)\T\#dEZf,K&H2I/6W(XMPO)[6bAYD4\eSe^A2XP)eSIG=/dd8#-S1+\RaMf?@
ZVCPG[Zg3CH6AUC(9;6F4IP66X[A8#NFB96ZKF)2+b6ED\B<Mg2K4O#.BPL9LS#O
f8RC##eK.;YOZC=(DK@.H,DMf?MW9VE2c1:@O+?^3E)G=PR]L?1f3S?(F(@JQ>N9
4^gCHf\X/M>Ef/Y9K[>XHbXg>e<ASCSQVS^U8.JBL.^]N)bfbN7YS>bP/E#7Lcb+
:UTK\TP3><Zf2/eR,@7PJRe<-aE3WYJc#F5U18f.(=[JF:QbC85LSE1aLH2Z=;DC
d?K/TQ:.g8a9^62;,C?+V/#@)W_:R800K-VF6UT1L:bGSGSM\aPcOgOD#K4=XA7(
K1J)]D1V,_;XDK:&FJgQ_/3N1-9#6)Eeb:Q8GCOTFPcAI855H>N@B>@E-eJ/7F+8
Q+N1eMS@b7E2H2G7K:J&<-=WePb46HV@P?S6,C[<)4OBO>;VF3,2gYZLXBfNg:NP
g@2[bHg>4Q7S=KEK&b7(VfNf.V6HZL)PL-EXe1_/FVX0/a:219f6FC?X9cA-KWgW
4)1\NGJ6@<_S8HFKEINP43BfOFgZE7(bAJ+4;T&,9UKCU@GAI_A4HgdeH^F3O2U4
(Q+/H57NSGOZ]A@1^gF=L&0)658SXL9^>d0NEb]6a2YGR1IKM;#;=D]04X@F7-:Q
=;5YSJb5fL)C##d)J]6Ub;;I]UJA1fS=O6A73D9JV2aU4:/;)M+9Z5=>/@9HVN7S
I]eR^PN47H38YeKaZO3H[b.g^];0f;:cTI012ERFTF<TaL6X^4K]CS^H-0-86d=X
bc+Oac@XPO-WTJFgMM-Bg\F;Q_Z4T]T+TG^G<SM\N&GBKB(8S^JPMSE?a4+-NG:C
G/NBePg\b5:W#@ad1VaVPX1O7P2D2UV5dZOS?:7-X]H@C0<Z:#B+e,Ad?J[#^(2?
/>R6fgWUg&8E^).GIJ6X[GS)4D894Q_<M)W7]Ab?eV.X/,-K^U1.2FVdPbF=:]Mg
GY6<-2A+dA<c;WQ[C^>,Pf-\[-&BTF(2>&RgO[R7J-(VJFUaeg<77UDU#9<Q40XA
MKA-84939a6g(]Hf6>KAPeVNaX#.NE](aaD5eOec3.PD&T&8c8\\;:HA\ERb?T/O
G[B7W+96,#SKL&_^D7DO/)&,_V8([Ife4U^2>Q072>@4@42@f:DCKfc;#XeB2:9C
M+a2SMJW_PYZ3);SET#\&\Ce[CU/Z+H5@#Y^Cdf5S2_Y:^IcH#T-TL)\g7HP3-bZ
PT;N0L<:)X.I:3P+X.C\@<U1\?a[<Fa;.7/U.Kd9ISF>30gF1PBF3b9Z;?L<T=LM
?\DdQaBeP1,2NLSNX0VKMgXeB.3U>+:W)@=MS+\Xc1+[Y\QD4KAb)f.>5XM8\[T(
VQ0,M:eSCD-^B[c_Mc+S3^Ng)HU2745W7d:JFQ2KeLV36&YA@]((Z414Lf.Y6\DV
?>#0<NYKR)HWc\[b@&^Aa^Y9Rc<PB@R7GC,\9,4M6U6O.=\M=4+HbP4;YI.g4C4T
=c\6O-L_0&b;fcT]+XUGW?&:O#FXd@=7@B?3WEf,<GT6A7?T?a.ab-W+G\G)b)(L
QV=4N7IeVd#BMBdTK#GLL4F49#X1HaI7BF-,H\\Z+d,c8;)^f?7FgB/79gE/-7WF
R1W+fQZb\F80?Z.@VW#:XDf_9;N2/a)gT7VEUVO+Y>N6#UZ8VWPWd3b0])J)8S,)
f3O83:P?9.77A#e?,4&_.g=PaZDCe?A=d@&MD/<CEIdg@KO-]@/b.WB(Y#L2@#1T
(2><6:N@ML[@EFdg?BMXUU[XgWQ)1KWT9dR2Tg6g13QYdLP@SO>g\.bcO,g)c/M_
6C(GW)6=1_GU[7a@86Ca#FK8H:K/7W4/Eb6(^dP2BY+]S(5+8f_:SaFCMNd[KTL<
F?JW=<c6@E_(7fODS?(?K6^eW+8OU&XMg&S<Y<[@@2O@1DG@/#<EM>24>9IAd:6R
)SW?9J@5geIQLQd>af6IS?OS[.UBRdZTN<?;9V.KOW\IQ9D>#.FAa:97g:_<-&QH
X7\,@0C:RPT=QV<6F#)_QSMU@UTW+EcD8@R]RFKR&\/C?XE9Vd(8)&^75;NeX2NU
\WbNNR5WfQf6^W^+/LMPUd5XJ>W;Ee7]_H-1.^?A..,N()7T:-VMQH9CIWb0:H1+
)=B@/TWM+.L3+TJ8ZTU8g\fN81[dfg,DTfNTbR\AfNMSB,;2@=eeWDc1P1F/2;6F
S:LMY=QKPFJKYQKTY>/HO_1:#K/RZ67dcAJQ\C]gM[:2IA33WDPZ]8@+Q13-<EHY
\<9\9\[99;I<AWce=^4<1Z]<CWO&CEO(B?O[6->9666f:[U\BIWHB1^5>:X>_c,C
M8#>&\Hb=?YDe(R@1OX88c?KU2&/Y_<82ZYO&/f<W<[S-][T]S0ca,C/AOS<4@\)
3EbCML7&>W72?J<f#0XNTe.?;A_d,WNE[KQ5UO/;A-L(CM,2gB3E1[/[&Q#/3J\R
76+I+g(+LeGJZ1g^N#&dT5\UV=Z7fCFVeXAI(N)]4+T(GV\4S&,dX[@E#7X5G,KO
f;^Q(QPR171^@7@Od/\ARD_[a+?cUQbe4MF@BL)d.]MSTM?6U5D=7GUQI[cGTXd\
QR-a+b7#e]Hf4U;K=Bc&Z1g2G5\A]T/Ca^bB6P8?FO)ZS.4@HcC)Nc)ZBP+-A27@
TZQ\C7K6U52K/3Q(VIb#CB:A;8&85a0[)A55>ITR)=+(T#1SbW(L/e<_BUa&SYZE
P8U.GSZR0gU#.:.BFeWRfR,S3>8Z(_Lc^NfJ)+0/@,<FZ.6^^&TEOGN\O[-KRBXL
^=R?++]N3:5C;6JTc3TZ7&BU1+4,3gFK4ae>3B_:F4<H<]^)6(cPBV\8Xe#>+2g+
e(bC=a?J<SXbTHF/A,KbgIWR_&^HUB\ZAPa]Y(JF?A#H&dUMe.+3RWR?eR9:;E;I
IAIMXNY^C-MD\H:5cg@>9LE19>F43]:)d1]K)1)b4>619IG5]ACcM((MZdVO8&/(
LR&af4_>[NGO+\R.&<];.>Z]0@/#\IDB4[H?dV(<N5Oc:Qe9A_,1F<Q;DAOI&\(C
MSRb\=KTYRWQQB\A&\CWC82,4+KB>gC=MAabD&b]0N+(;1X;b(,E9YET-Pb?]Fd.
8dODfg6/bTMdEIT/X&WTR]cLc<QQb1LHG)?6MEHZ:=4NT67B_G;Rab61\a5W3AeB
;EYe]S8L315H,M^-^\C2UAZ.RB0A]g9cY/eI]ZUYIG\H5P00#5P?^=RM./VN,gHT
B[?QD,0(S>LIXO0):7Bc+<H7?D#e5eK:H6GQO?-W]IgPUUEf,gFALR0f,NKL_CL-
ATNJ<<b^H/UXJ)ZLHD0:_b,EJ-d)?MN-?<=#1L+1&8DK\NZIM/\]-H[M;W7A3Q2G
N[eN30?<fSL^YZL#6GA?_T;&:?VRLO#S7e_VLf-e3[K>FPc,P8H3-<bL7KKfY;@&
bR]d(JXb9dT]5KQa4A_H57SNH(M:]H&[+0bP]SO)MV5M6,10e1@UY^@KbeTa7[EL
:U(=XYUI5N4C3GfDb0;e/<1aC7/AEN0P#/BSCKMA3B+gOJcFG]OAa@J\;DaF/6,O
:5\JPQ07^AB;ROFM2YJ7B7,V?P#EA6(25^<I)ZggK-9>+a-[(>?[=dfQ^)]QZb/7
V\fb-Zd.caTOGgEJV.N9WdG1<be4EU+bEP?W+bYC,)+R/1@2J&DO?8:7cg216cHE
HbG6DbL><Z/N_+U+<>]0PT?aA^/,Yb8R77C_g83G\TBdKe]?;a#CVLc:@[>;YM]E
;NgGY3C;YJ1=0]YCaFFPN@7F@Pf.<L7gRR3bMV^(V&FRL7N0FBO\5Zfa])<VP6\^
S71DZJ_P8#A8<9F@MS-U<[c=BNN((Gd?6CO;.@T>J6)V]0C<P#]ZIJ@1>gSHK</&
.BU#5PUM[^P-H6Vb;D:EKf.#885EG79@RdO1g]K[[PX/Sd\0N>a5cKHQYMA&;&g<
@O,c3F<OXI@/fB#:9PSNOAFIdOaRf/QL/^.NUDFcPE6a&NPJ=^N32<FA25-O6R\3
^6J#bda&WK^ad/HWY]7_OC:PBP>B,,X#O#:T&e>[J/:4+DOUM0WD#EJ^+6,(S(b(
]C_V(G0#c_C.X1#T0_NC-g6QX&1JHacXEXA)0B-P2RaA6K]R5H@b,fCR1WX:UGS)
W(EY2R)__YZd,LP\<.^ESI[O5=gCYa.>#AL?2G5DA(Z..Q:Z@32(>?H>7SV^)A8<
FB-H#D&:@,#NfLQJFI3?1WW9=PBI(JFTXKdR1\fO+TX?9c;)bI13<^7_g>3U8cHb
:H&<AZ?Z+U97C=M#/A6;D3(&QZMEQR_^3#:9J/Y,?;dXMV3W.(C/c.b?,R,MN2;O
7ZIMP\\:BPUeeJ<eA?fMN],T;@791A_0V3O<=PF\PF??+6;<=Gc-GZ6.C6eZ)8[;
FbQI3;K4)G&:_O&NCAO23I6./.<Wd@Z5?30&KOEggLT>Z.2GJT1&&0R3_<NL6Ef0
>UD)[\8I]#H[8+e:Q+8AZ][V:8M@g_f;2J#L>([aST4Z3BIVU:[g\CTgZZ:9Y8A7
<S\Dc=/YQIYX97I-d=OUcf)P<YdA)4JJKEC&76IF4XOfWVaG\.H7\N3F1>H\I@SZ
?dP#WM<,SJ]4>5:N5a;]D+/_3_,#4E2QUeXZ=eE,QS@(W0PPfY4=Z)Z[d8Gg\[AX
T#UWV9O2cOdEW?aY:^KZ.6MDAQA5\DDT0<7:PE,e)Aa./OQ13bad_JE<Oc=,XgJ0
O>@U&>Y86-09_;0JEG)KMRgQ-0HCI:cQN0/5YM:V<^H]:\+<5M5YZ81CUT\RMF),
;UWP2RcGH=NTf)GdQ&;;?^OS+2N/8^];THU=Z.52[SCYAAGCc>729PL<PHX-26P+
2A+Q(SgU73df1+S]O^O-YAbZ+JQJ47H0d.bdaTUGL0AO>C@KE&>>.CNJ#a&4_D2;
N_&1@?K9\7SL[(VP>W4_R2Y:daaB;Ig=K;2>-P:=[=_<f,GKAW[(])/ML])47e1E
A6eW^M4IcWb@.0Cf&DY]PN]fL63L0+]a\;4T:/:B&_,N6H/615CWDGRM[6WIA]P7
E69PZ8Y_-C)MC5EO-:VfZ&=0^e.7\(bIZ6V67FO9O&PG_DNJc8W\)H1cEOdeL+EC
cDV)&E8QJ8Bfg)EDOOAZHO/fS;eF=<gAe/#1^@/<[;HfU89ALK3>d]:9YE)c0-9J
<_2.IdE@],Q@F34ZUQS2Z-(W2dJOBHLE;+caN0E2>WXa[W]NBF2^0#1KN7:df:WO
ceSM)gYKE^[HNMSS+AU@/+OFZ\a+:\1?1Z3PWcge3b:DF;.F=a1GLNSMW8I)I>[N
dXG_D-EW2d>]SPM&3Kf^0R>E>afUQC+9U8a=b?Dgc8H7+K8\S7REV:]_@-FSMfLN
_31VMG,#@9D1<c];&F8e.C>-SgSdeHH&;d;eB7[9UDKK71HFB=OE;3/Z2E<D02b&
NPPVVgD/8:C4YAa];&Cb7AQ9#++>PB1Hf2/:BSc<Y(YY-I4ZVZa(74W\FFa>f21B
[Q2a?NA3F3ZG3/64:#W1ZaQ/2f<]M.KLf=@G>@(-CC<.?e<G;P9WS_999D&ZK-]Z
DJ1ZWH<dO(S0F:eYD4NeZbRbfHfcdfEL#=>/e<0Fd[(@FIP:a3A@5^CNTGQ8\,/4
GB?Q-UHHTJ:d:C=H63&<Z9V^A).A1C,H?5G?+a-Q_1FDI<6\68<,=DTPf^ED5:B4
&@1-N]+L>LMCKWV#WTaI-DN9eaH\>)J3M9Fe@?fGYOG-1/J@8PK)ZKGFF9gBb:[U
536L=G]-D]S96X?P8(L<\N\8T;)IR+SUP8CS<g.b)7#]Z+;)+Y?Z\=&[CKdI-^L6
^14eMaX7ITW;dFQOC5F:@JAD7R36?=3b2XD?QKC5_\_R+3G6CR3fT_KK1)3&:W5L
D@[\3(<MN]/Ud00@)\b([,P(gAGR/]W5\G7F+.://G\A]#(\,9_Ga.GW2_DH_7KZ
E17#?6QP[O\e1YO9GWQgR6&9afJL0?.&>1Ied:f4T,=Gg]2]<)\Y#1/#L.Mba>@F
I>WF4>dDP8\Y0&@+B9fR(eO+@5S:gOKd<-C9,>>8A99O.O-RUeW)F,#JUKZ)<2Sa
b1CB@.ge9cS.9g(d9NH8(?A5+BV?eA4(62FO&BW8eIEV[c58,ST13MM\2/V;I?)P
-dMO@#Z;Y2QgDJ@=SPU>7GWFC=cXdbO6gHCdBV0V\SIH/+_/NN8G;X#3?H4-/N[E
L:.57VOO;]?+e_S7gaC[0I5I;_,IXeB/Sb[S1QOFBd]6.@Z)BZ+FMPUX3Y(TZLdU
G>=#0G#gNAHdMUBF<e]e5.,RBEP&O@PVWXL3?QA92M]+CMM3W10UcSg7HcebQ<_B
-dA_Y_-Fg9EE,_4HR<4P9BNSg,CHPE]LC+.5H]?JCE.e]:[(DNPV5bTeHc)Y588g
fa;?DEba]Qe<&.#YEU8=:80:LT>1C,a(X3d,/35c:;+DPbP2ZKKW:G0G-B]6X5+9
;IJ#-IYBX/7?Yb)X2(A]]DG.A^,@DTKf)d7;0/3<&F;CZd=dePUJTI.,B0)Q7,RN
=.C0/3Z;ccH#6c\AXCTEefMRF]2R0>W1F(<T_\R@+Q=g=P0PG\+eVV[caS9d:O>b
E6a7\=)bg;(+U;Q:;[[<Mf5_bMBW&>@[E#8?fI9O/]Q[3_b:E_4(QC6BE^WDR;YM
UOIGDF#d/HZ.SA(8^>N\,CEA6e7>a?89R_.AT2Xe9K7D,:9T3Ue4eWZ[cZ;AA:WF
)ADFH32:_#,&DBZRZB>61D;]9@.Q,GR9H9H2PP]W0X]OeQ6JBA^<P\>5XP^WT=KT
4+e>UKI+?D&S&Agd3J_aQA7C#>_.,04-BZUNS237S>X@H@.J@_A)U5e04Y1e--/(
ZM>Q9=RO9BL3,e@gE@#,C\#M(^+UE^O9E,:N]L8bUCVAZNCW47>U\^1.)S6CUdgd
d@\/)UaMT_^Q/C3+,E[IS?0:^T.7eL^4,+2UZENIbMV\&O)K//aA/5AE]5.<4;9c
JgLV8-Y:CeN]NSe)XSGF@7,5XTSc7J/4;&+4WO_(0d(4/6.0.#2Y#4>bM-YX_d;6
8OC<d@.2^,^2N0<59+V-5HDfJ5g/f9MXN^2Q3O_J1B<\0MNVZO:@&Ia]QAJF7-?D
+8#)T/:ZM0KM,V;.=S7?2_3NAG6<5VH]W-1&OC4EKIA4f44bC&UAf_[C]a?WG_Vb
PNU2@T0?C>OXf2.a^K6egKV[QBe&XCd].2EX-FGZV4#]7-D,.SNXd=A91V]A<[X(
WaJ=IR\,@E@aCXUQeWNP@dYA6(/R7bN8#(2ee3a?/8M\>a6ZLTOdWfB.3^#\f^<9
bAWY5.HbG\F),3YZO7:I9aXM\]QCL:0Ae3?\GGB5?9-(=Od@HM8_(ONeO?EAG>BS
4K1-H89_WF6G9RDHHF+Eg44RZUT.SOMH.VdV+8K?RE5Y@>-<;+9fbS1E905Z:XID
9@?H<AO1P-SET/T)b6UcdELEXgY1f=d.JA0;&g-/:GaH/+B;@SVYf3ROR1EYK32G
VPH45^+T(17?.Le=02PNN.88f]K,XC@+BE<b;aL_O-<_d^WNa([c2/\dB=7I.7c+
Cb@/]Kf>[#3]B4BQ=#UBTR1Z4?^6]Y6&^RZ]S),LJaf0d<T,V+#+DN(;^=;\a+Ld
AZ+Me3<DF7eSNX?98<FDT(+g<3E&2SA3&gNV>>5W+NcVFGBAR]]\>Wd;<9Gbf=ME
beeZ8\@6N+2@:<=_e<?F,_TGebDN2@IRT]a)H-2HHP@PaK\_?NKONN/_UN7/g<S/
<eQa,Q;AAC;[+A[;58.0(dKCD,,2PIbP-XF]_gAW_7YXGJZ9[#,/ZgQNO6\]@GUB
6^60?b=.L5J5SEP7:L#&FYQ^G5&YG?D1)9?;3C^0K<2]FVCQ+X)0>A#ZaLW,^LW,
2=cIVNcH@KN-(QXIJ[>[[1LL93IcS?/(aK>T0Q?RR_#P3c?VX:fE:ECX]];a>cb>
?PH^A&=Cb&_S;?(0=:8N]?PIDWH9<9>f]2#?QSDR^@9329aB(&?2X\O7GEV>:fgL
Vg4QD,D]ZEKV;#BB+6UDY_3bM61eQKM\YS7dL/bSH@d44#V4G9(aQU#\aUC#W724
8[6FK71HQ\8eX^+[Y-Z885M31FG>T>@Y[DJ49IXPabd^\YSNVf#[dNMG+62E<8H^
OYR#0/RB@H.Tf5CJF6[KW];L#&4-9d+[Lg->EC3H;C.eT=H,ZJE#b41T:cE=f(</
#)(T0eW+S/.;-MIOR:\11gd?+&04]+Le)0>cd#NCf3I21U-6-A:UdPd<,aAIM>?#
.a\@ZY3Q#=LYU>X=Z?L]C?)g>0Z98E;f6?&WDNf_ZS50)&,N?++:Z\PU(e@Q516-
Q)0#bQA3QR9D5]fL83E\0E5Idg;F2GYR#NE0BQ_=/G(UL<SZ2YF)3^R5@D>F#Wf_
+=CIIZD[+J=9R7gV_:OHNX3BMd/ELV9J21YV&DU_G3<We3bY#W4]@-#[KIV9+fY2
VM492bH@#@feM]22RP3J>6ANOa@&_Ff(g,)gXLg381<VDQRY\f]&1-1bF=Dd;C&d
]5487d]^;R\D;8QR5UJ(K(GF01/d]J_54&)=f7Nf[eQ;8^>>:P1\Wf8T6TB?OOQ@
H=^[a8>N[/L?ZbB6AX[LD+TbD1GK_GWP9@Eg-[(I=(Yd99DOI3[N5F)+b0@)d0HR
PWM<+baRJS3^SQONIaB])1U3ca\N).?A@]7D4YP#@9X_FIYbEafI^f>T-[S@5VUY
e52I<U(a@XS[4;FeSc7Id(ag5QOJUfP:d<A1^_[2Q)]OLf4,NJ^caR4KZL98IV:G
\U2NW4Z7&FH+N-X5B.K9M\CQZbCGKba:@VQ5b[>DKFBg_&(&6c[5C(,=A0/Icc&_
Q<fJ:a)_YRcfXP=@^^@U::3W^+1EKdKM&^<I)X6-Q7<ad5QSPE.1>ED]I--RV,eB
UdgX<6ADDGb5U]6&gFJ24MN2&5gJ&\9\O1a11<5D<MCINUSW^[7B8@a^_WC&GY4K
@(LK-/e&=Z.fZAG0.2R[X.^.dVK>b<Q,CYg0e7Y<F3#Y@9c&0>/3DTD50PgX\?C6
g?^f[EeaeQ2IfDA9LbKQ)Z[80aSUf#9IZcV@gDKHc2OQ]MG:W);AGXFE)3>^+7.4
KZWP_cP0Q(Z#=<MCd5-(^4MA3]KV=+7W+=^,;G8W]@R5+(>7DKO(Md8Z1,D=@KUW
[RE&D44<G#)Y<ZUO8-Z1+,LGSIA<>KA4aY0Q+UM?Z0E.-c).McI>FgO?4E-)UF+U
;0U]=KUe;XP2K,(P/aM1=6HPKG.LIYSGP:T<2/5RD(IT1:+LDR2Z?RKG#I<;#Wb2
_dR(L-K546>@(-^ILVbGRK0#40Ba\:f2?5D3&3FW\[1/?2A)LD9CJTc^QD#Yeb2Z
>B[Z=M[7c>5<QQf(-g2KQ3a[Gb]a70BGe9G-P;]V&#B[.&;&^/I=.0E_##bD?V))
aA1XOJBR.H\3:BMa_HIR3bNg+M-K4d/I13Id22>AZ[8]8++7WSUN;?Ka-7\9.bU_
g7H,EIA_>e-gI<#80&-OM<FK9aCWNI7;#8WV\/OOU+U0a,d+H0+JgT.&4AL;f;_Z
80+X.,c.W+K<\cY#C0><ST>J1D&OR@QA8^DP6G(YG.JEO=CT@MIW8E3&(a<(5N8f
\1<49P6X?c9MX7P73QMe0cJRd_O/6Hea3U9eC)/3,Fc>,dN172bIKd8;/JEY7SFL
5J(c=X?TT.,dG3G?aTM1A?()K@d(8.\e(ZgE]QLLDRLJ3<ZZK[PB_RQ,bO7+-/0^
F>^19&Z0)SdcORC7#>.Sc2UK=H>>-TQ\AJ3#-53/g=[ZZS)A27-Mad)6FMX/0JAT
,3Bc#[1OWA)ZQ&RV-+QP6]cU)^B+/\>@ZL\dT736@aM2\-+[;PRP5(OQ.3a1d:fM
RQ-/1OB4+:(F(13Hd.]S_9#/4_Z2gM58N2gFaK-?-KJX]B(P[_XW8T2I5gAS>>3L
BOOOS-YD7F#]B_=a_=&FQa#35fV4#(@7\[]^5d_7N44RY(N)a,Se;0RS-@_Ca57P
1MS;1/0+PE&IHK?f\\?GAD?@2OHXHe<11@2?-9EPTY)RaN;2O(8ER((HURLL<U4,
SKEJ&dEcYH&(25XXgbeg82H7e#CB5.JRgPVLF^WS.5IJ2Y^8Cc.,HKOGgI3TUS]@
QI[&6=e@]U20R-7D-R#d3#OO)_;.e7Re(gD9>[(&U)aUCA0378\bF]\5^CD)L&b>
&Z1F>WYcATJ/>;V&b6C(0(.45LFCbCe8S#613ZV6fGJP,cPRAL\VB>-KQHD;TIT4
W1gK,LBKHPF\P&VW^3U;S]0NP:S\Q>L?[e-+-_[-3FgOL)FBA_<U=2CMd&8#41>g
/-eH\^6gML_<-GQ2+_F,5KHJ5<MQM<gLgg-WERW&Eeb5UN<3(1R9a;3).8XHU+F3
IP4g6D8cVJ77&&.\98Lb+e9DO]Z&F[,-C7KZWX@T/0)B_c.M2R>S_fMJ]ZV+@MaB
f1-1[7KR.aJ1\_5PSUGUPVX-SaJ/.?[9XOSQBC-Z5^TLM=H1ZY8L\CK=6CbbJeS4
HO_P.&8,8/-5]Y+Q_RHZNSPN(CK]J[NDV_T?GS4_A=+IE2)=d0KLO](+A/:M8C(f
X06JF=@;K9bFf[Yd;Ra>0O+fN#IT4<I(H;Ud/g/\W<X:f:df3fONbU;L]+QN2FM+
6@c#LXAI_W2GMb_6+?7(I),+8;M#]QaTT.3b_KQ;2^SE=B1,aW9W_ZJ:B\Q:_Z.<
/7fW015E\d0d^WR+N?)^D.J1J+f0,Qf=QTH3SI[X@->)E4..W3U)4W.?fg:;3SSa
(\06BCTH]W?62LFCbHOMCU4O7?QL7G00]JEUEXLO_8>C_559g8?\(WLB@P\CP#aQ
:gb0SGeQc#\).J<(@dZ6FZ^ObG]W[7F[=<PY=IV=X-[<OJC+A_Z8+McJ)ATBfK]I
U<TNcR33O;UI9ZL2?5B-?4Z#LO_/<VAXLg-2D<-&:@P?+Z9RAFZA(EA&F&D;R7[3
Wf;fY1YQ0]L]CLQ2Ia^Z)Q<X7FIHa,If8f1?E+e,_D?)]+fQ@3b_9L8BBT+>6H40
bD74WdA-)f2a4,Mg&/c+@.5V_Y\)GRIK:+?f:4:LPM)b2EIU/9)&D(&FL@2_BL9+
@J0;4@NB,^F:IJ0I+2V,Z2[8EL>?)=X8>g(MQ1ZE>2-5ZJW79bAZ<_RVTW\.K25(
QIQ6#gC]Oa(#E:\X.eKU]9F@W&K;Z>JZE>_C@E^e1<_^?E9:Ug3S8bbMYH9EOXf2
I;6fAWG138\A5&?/K2@-;?HKJB/<0SOM7)G=[(W,#[M<b-2.X1ZgX7U3Ad=R2+.1
-ZVHBWR1@-I<\c>B3[e:QMIa>IB,+BX0DRf3<?+U>ZHZK=X[c(]COeN)B1MU0Q[Z
9EXeFY:7?g#:gb3G[Z&eK5g(U]Q,#1e^J+gZ42\<)KN&I/[+[QAEWC/eZI9TV\N1
5Z;I966-X:NU#QPK>CTL1eXaS3WU@:6>-UWce.<X/CP0\32a4TI.aFcP_Q/ENaLA
G>,>E9SV-NJe8#O,B;+(FH?E1VO^U.BKW2-\O]f&F</ag]?;.A:28=Pd9&YYAIQY
2W?2YS:A&7NJ8(+@H?6dT4_E.7D7?T,W1Z5=gV\,ML9K]TIS4_TD1.SV(_@83f)0
T/7#_-TV5^:f[KgagU6.;9dLJDO@T,;/ZN:R<(=7DX<cNF4/<X.JGB(/YX(^,DTb
&YTU>+=85d\V]I4U73E+R#>\Sa&1O(FR)O<OQ&2P]&L_:c7?J7IAU-Y6,5=KdbUE
HbQ&\W_L,:(?XC=LbeQ0]G4Qa\dL?^&Nfd]<1)fb<W?UP?^P@3Q(,:ELY56;bU?]
MVg:=]A[WKG8\?^<4&DQ4C.H.#1FdU[#J->/9IAS)C;6ffC?O/&#9O+>c@SDgXKb
\+KH:X&XF,P-;ge5J@H1d4&/fd7_>P.e(#M?#;-@M]T+?;.&G+a/>[,G&X[6&f?&
A]1bZ:;_T@&5@T+BgEcIgTUc)b>8TaP@O_1>22X=-SfFI/L^ONS?I=g@[[cJL0cc
\PcdHJZc;[RE^WTPN[B@+8WT/g,CC^gbW#d?NZ\O>T77Y\W^TB;>Nd)3QR,Wa.VR
-_76S+R\fRZJJJN4b7U4A7Kf_Z?Kd.]+45KWU-M:/b2P8b/9#XBdg^/Z3-I=C-AP
@OdF&BITONeWc8P/Jd/NO;]-T-Q1E&/5<a01A_gBSI]MS0C7CK-)LQQ@e0fWB@fT
@:cfU1W=W#H-Z^U^0bG7NNO0MbY5-dPZK@OFcWIQbRVTE,L/+YE7C>6U9faETCQY
QeF[8:_1#d<S_<e1:CRVJ9YC&>S4cf(6>V[U54SKVgGN0Kcg=5Q))Z4?>ag)G?CD
&E8/&7Yf6WQP<5(5EM@,5\G^#G&F7@.E;5?ZZd[E?91U6>Y3HO,>5.=V+Sf#WUQW
3W)TR+9[dN^IEN^F;WW1VYVZ[53FEDWB(66O)CW1^0@T/QW2TC.?K_+a/5;W[.g1
HHD/T__+(bGPdV5LWP\e)Zg1675-^V6ET.EIK48V8=98eW4B.-C#<K>A:W0UTK5=
PK;WG.WX@+ZT\MN4RL[,E7X>=V>?(#@a9^[P9EKBAF/>)R_\_J[FQC-.<I1:6;ZC
4V:0Z33M\Y4-JQ_HYc+WEZ<Ed[Z(Z3.caXYU7d7X9/9Hc52Ja)N[Q^c>f#+E+baI
#cGCM)(:(H/T;/)bX54GBJ<J2(F3T6cX&_##HL9I>6[S.I\5Xc<Hb(WF1?.3bc[M
3=,,a?J33?/6E(KG(LJfK(N/^:E&H5b3dFE7N=FZ\F>gU)fP3D?=aRY2L\-fFM(.
R953d+A@9^ScWb(H0T(R.8<,)V>C3cQXfQR./N(]<F)2e+D>8N91-24A6(6:fXI?
:M?1SWQ]C9^OF2B3=#L98;[M)V(IDR#F^J<1VYZRKUT3Y3L;(U(0c>fNXU86FJ85
?9b<:&?HL,,a&1E>dE@aRPaL;dHDb43f4DRB-MIEg+)(DFL2XMM@(Ud_Z8-28;LC
f(?FW@_C/=@]WV#^,aCL^PgGZPfCAc3\ZY_8(R[EC?NMZgW^2HUUEGB(;+[<@?81
>,cUE>6b04A1S.KPgL7+Z1#VN>P_\HgB4R1P/6P-.]IO])EUE5>_TgUP;UaYQE#L
H@PQJgT4M,IU(+]<E;.2WQ&8Z1P1K^H##7SN5JSM+D4FD\3PR:\-4KJ@E/KW7A4\
(a-Y;2P.eL;-#</65a=UMKf;5CLJf+XeRT4#L,P(@OIJIK(3g+/6ZB5A24g:#ZDJ
65K8D4M7JOd5,KE+S\R4f42EKFOT_:F:Kf[Q;aa=9\_W87a=,QO_C5AZ.:N)QVPF
SH0daHW(RAV0Ha8S:2X@:e6L@\gU<I_P_J7//0:#72C6.H9-H<05[AW<[4Q>Y.6#
\)b6B3AIFHVL]^L#GT?B+7<_d]<IJc(GO=BOR3700,Y&Q03^N:1cD97LG4(=fa4V
S]=aHO>YM656UQ]E03)H;M>C&c,EOe+>G?N(fH^1:L4>g92X025dXLY7&EMZ4U[?
Zc<5e+?IF(1_87&2]>2F34A7++5MX>HT[LUG=dT1,:QT-EbS7FbaL8&,+ZbU5EMM
b.EBX+Te(g]COcY?^@SI8\U]4:=S?^E\\]+FJ79?86&<O]9Y&TH_fFMN9Y,J<FG[
NI#SB4WN7YCW(&V<0##Dc2J(d\@>;)K-g)#/84D:HbV?bb).+SPdUS;#VbU-c09+
P;YMVJ^;ZL;#AU@cfZ4J@3VNb,)?4)V833IESeANRg2GdK&,C]CWME7fN&OE5gT8
QMV8.@JQ@KK?Zg<+BK2PWSdPd&:5U6G3I76DL3#81>&.OZ;MD5^PZH)2U#1]&7ZA
PH5NVQGc-,a80b[DOT2-&JMZRc&H53BX,1(B,e)3+1IbG7f.K^]f87N==S=A.XPc
:f^T1(2Z,7H_H@KWYHM4WPa89?74&)#>=6?ZKB+&[T24)A,-=<)A2<dVL4SJ+FS+
7+W>@,gg@dB(11W(RU&QG+P819NGTV_P==,1W-YbI[02T0]8PIA]0(9&&YOd:\3>
0GCg:0Q?J)0]/X7gUU]@]^UJ-@F/.&dbUXLM/]@S[@GVMC6O&_dS4\1bB#TJ,Yc#
&ReFP5IF;C5/W>M)bQT),^&#>LWcP+;53L-_3@AP./]BIWV=]0]_,CdL-:b24e\-
c):X57c;XNM.E7a],C@FCUUaAZaT0#<;bW^b[#<DEEe:,>UG:5C^SNMUA2JY)BQS
fPJJQfRQB6B-RD(<3c/]g<aEG;N?KDJa0TeA/d9L\VZ_1IV&)+cdY,@[0UCF4(AC
b6[?TS10,U1.BIB1bZ.KPK=N)3cXNgd\9Q15TDI3g8Y:2V4;[-MBHf3WdgT,(2IU
1J[f\V^/G(4^dg64B\2O[&#4VLMT8GdcVfDULON.ggRYCWBX]G4+07)g,O/e.G;B
<];X:T4QSQG7@/B.K[b&efcfQZ+Ed?#&d\4KF>LMJ<;K8CPE^U_K:6#Rd&GPUY_g
,-\@dV1,O?-=0@b=3>6F##D^EY&X9BV-#0)B1V1dYJ,AOc0H](46CIaP6=;;e0J=
J[QH0cW>^NUGEN2(R1/HE0cKLI1_#BXF;MRLYRS6dWP_9QXFS.ZMVIZ_H?Z[f(6X
2C4M&aAMb7N6W&(GXN>E;/.Y[/VP<KX>X;H&7OAV^=HM+0L0f,]e#.]XaD)?I;Df
9[g:4X,M&+.;SRSI@+cEIfOX?D-e9^3HS+0ELeNcBGbW8bJUR7N2BD-?c&eSM?Z2
BB]I/eBY3XG5>B077>+9/ScLGSN,#^[5B-.GJ6Ne5GNPJ>Y&+Q#^FS8Z)==AZ>=X
VREa+B7=PEW=H2gN6YE@.NS__ZH:6#b4&c+W#]0,f.V09V03)0B7Z(ROK9?g\Ug<
H]3bHV;KMd(dVcWY0:-]SMR1.IO^BIeBG](KKI<M1P&,C53J8gF,R,N/Q<Qc3(LW
G3;]OT>/_SMCZ]<^9e2cd]@P:1N^f]\YOD_BB(d0=QD,?U]0>+R:b,f>WA9TfdMB
K-3L>b5BRa#WQ?9=bF(<FRX7[51;4K1U=+fX#>.>QX9:/B/&0M4LDRH/5ggf1+M.
Pc\)Y3DPF/C0.bQ.e)^9GR52K48B+[dIN0f-L,X2,F3[EZc8Dc0(F45e/,BOf[@X
D).:GPIKa&]9d[G(M8G<L_2(5AJ?g6/e+)2\H<-IQ8F8g9V\:_0PIR1cBZD;,GA]
?T#N[<_TV+J:>&1[WM<[f2EE/TMLeK36UeGI]RDda2HS.&LV._4AB.dDRaU7b).M
N#W-\VgS[cVG>g^[3)F,1UO<08_6=VO/f0;OI5H1]U5YE-2^a1(Ea/MCF50_^WgC
Cccg4/=[aB5_;YC#MUcg2@O@:+W(<6>K(UIPX@-((12aR/68fS7AE[e&>?Q#M<8)
O96SJW;E2-EM@D5<T,MLQ_Q4@L@5^[[bc^KfJ6SD]YPF(65VNB\c@Y?HL9B+(dcW
WOBZRHW1TY1B^<U>I+=>[>G)IKbFV_>M\/J4CSWMff2,M9\gbSF@;5/A3H^\;AY\
JUbWf(K=SHF-&MTR-]^B,K2]-QOc/WgDNWOc4g@FP[T+H/Y.F[5gL#OK[ZTJO\b4
,FH@SfC=DJ8W[-1De^&L+g?FI.>(#Y:]E/WVM<5)M<@Z5d/fOcfbAfT_3FA?4W[2
e?2\XN:36W^J9QPKYSA?Q:J(8E>DI@16I1M0:R#:+CF\APSfX4S1[;_VWHT;1FQ-
)e49H_G?dM[293_,M2[MRR]R[+9>8LZM0\([[__^M43&M;8TJ84UU+9@M5gI2.HC
AKCDLG1D)Ye6>]97PA9P-\K@JBd3Lb[.OaUY.0VH;=7f^[4B\4J>>4a-E8AYQ\A(
JI?6>,\61\&D#699WH;FNCPGab1\gDWDW74Z./K^6KG@2&&OIFQ?EQag[=E_ZUAR
,/F<eEe]ONVBb/2#&QGgA_JQ3/.D.C/U.#-I0SXMX/a&B<^+8>RWS5+UaQF@<E7F
W9O5]XVYTONGRg-HOeWPB>;FII,[0JY]OX3T=RRG1VR#LYVCVc6E3]1J\36R8Ce@
LV0<-3_OZM9>-U]VI#A^&/E8eE/E3&VbK_b[?,-?Fe#:I@&Ce\:;I3<5VY_2N^3R
7Y>@/OR7\NG09WM1?[B#,&;\S7_/e6b2<F/KGV4X0gI/Pf:[dHMYfU2A2P[OQ;^c
6UTJM9cZO5D3JCQ0_LG5V\/[>f<]:A+GW:G9\gYY1&5#:(Q6:ZL5#K;8,_\f&V4:
(B2Z/7d8,B[MUG9&,B/M0,<6P)9CV9C]XK_.E-W&ed3<N?WKK2AO>7Pd(Hc.;Y/F
8Z1b+bf5ST@AN[0<dK8\dgN7bO2+RE-M_0R7/PC41E51/=>OG#@/T\)-,NIe6e,C
2,R;Y9@#5.GXL:&f^._D@#+IcQ>@E8@e2[XMU)2\-,9Kg@;FH-+IH2OfH1_UN9,@
RFCCB^Y#SU5A5#?bTKN^0d_7FK#\UU#I),BdB^c(YVA1UG1d)SaF9gWFba8a\:V6
D\VP/Y9LVZWgMG[dH1[dF,<G8dF]UTT8)HgAMIL6>D5^\3_/I_JW5=OA#3RNT_Z&
[M+,F\c-#15E]86I;&AR2BbS]NVeDDSTIQ(ZM2?VIb=&gN^1K09+(BO?&3.J9)WF
K7)1#5J,I.f0>4XZA5=_DV9=WET=Ob:()Zg,=WRg+E=JddU>^5E7b_2K@0a^E4bI
WV6TR(0HZ@?4C)>.;XcJbE,D&H-IJY^D:8IcN\[b5EX2KcbcgLOWdfS:A03RD>93
L1+56[SYfX-H.C9Z^5ITbaCLcMIX#E<Z?>UGUR^cHGKSDb[M_T(5d[_[\114JIf3
WU.4V/@GCOFM(EK3FPI<b:&#:B8R7LY@B,V3)9[[YMeAJcSU68AfJVGS;W4ENLA,
H(M?Z]FcGe_Q,@591+LD:B1-)X<BI_RP&D@45,NWJ<33J;0#Bb)b;IV\TPD/a)fJ
c+:T.N2P]0MFYIHCI25c^WT6.R[QB^NJL1<Z=P.Zd0/dN>;K]38-:TD00C]HFaO;
:[<ZH0ecUIC5;7N8a?1dd^T4LRASDO.XEPe]]BdJBYN;W+#>(5>#.>A@GOO6?\Bf
Me.G)&X>R9-Ac=OLC[7S8?8[<-,-TLbFOV;]W,=@ee?7/HBB;H9Na5]S5(aQ1ZHX
O[N3#de0f=0;)ddg52EaOZ[5_P6RG//9[UACY9WF^1V,Q#Q-11T?5eWZgG[RH@WS
=7&_OU8VGS3++[QegI<T.de)X)#(FeWPK&F(G.7/XQ@+=Cgg[5a[L<>FIE4KT@3<
2LGgAa[F/7Le;Q-+:P[a2AG:20bdBbF2,)e,+GT76e:dWU7QC&\#aaRRE1&/UX[C
W#8-Cbg#H6,POTdYa5d-49A6/PQ<ff]#YN0EbN9XC]8([<a.@_-GGJ^]C/dK=06N
35[9?)c8BIU.>O3<\PF)EX)))U<XSA>YEL-1CVQNSI3VgV--]bW6Y@Og8S^M?0G;
99@7g;/O172VK6bN=J^e95\B3BZ#LT1c,.gHQd,+7NM:W_FG]NMT0^7Y]XPU#5:M
;=\LGVK,/DBd3]BXJ.,g\NQ_>,3O(#(3Ac/H1e4RSdASC=&M5AaJC,c?&C/TPbdT
[4FM^-gX,TO^>]NDJ?QKd&?,#/V_G)RgaB1gV-0<6:GG^KU0B>YFW.Q3]+70OZUV
C^QY7-)3VEU358Ud=.B>O]MLQ_2ccc\F5S6<_T?aFfg;K+:_Q@g\R,HW(f7+0ef,
P_ce45VVggJ]L^b+T^[V,21K>5d&=gWaI(B&4;[QOPa3,4?O;cg&>d,Jd4Db6fO)
S>ZfOT+B:b/FEAE[OU1XR]\3GN\FWV+NE9NFOg8KPIb\/0&8N6Ub,Z4cS\#SN?f#
U3XO_.^]L4bSH9[)34LH]:I]H5A-.R.Fe6)GZ2K8Z6EH,ZWY6YQ_b_2QcQe]F0[H
NBg0]72b<8GM5E4SA8]L8KLIX\0Xff6BXA[;?\E>c5>P5./_-,N0CIE9_0XIU/4M
-XDgQeX\U_6:S8BM_?,.17G8&C,g4PN.DNZ=-#M\gNZE+,:\O8]^E<TO[WNXgR<8
]J2Z8V-Uaf[bX0D:6]e,CHV\&YO@D14H<&-)QK[UBLX(]f;-O7)=>:@B+FP(O9LP
0?@<VEDUB8Gf\HHIVfN:O+09HE;\NP3d0gc+<c]Y>bI^;93)4P.UVK,1\GW:-4\1
U0eBNNKNVC?Ld;W=2:>IZ@OU]M;eVH,]M]=2Z)ec)D3>_aM:O+<\Gg.aab^8C<??
&,^100#2;b&O#H/PTO:7O/P5\WE;P/Dg>&d]LF9Z?:=N-F=FQ5N,&>MDAS0ZS2:0
aX@>bZ^>JUY?+])c.F2<L-<LR/))B(@@/)+VU6cFBgRBZW?]W@ZJcK;F,-8L6L^Q
^:T06@Y\6O2_?+\V#[WRb7:1ROb]K=Ld]OT[/cC8=R\SHL59W5;Q#JH@?CR4[WVG
^?.ZL&,YPaeafI].-@T1F/.;OYKg27ge\K_M3>&)aK==Ke9UW-/8_Bd0XTGB/=3T
SF5CPa=_18U0HYaP2<MKP44?&)O7NI,a/G<5IG[O_#^W@P5),gHQWTN/)K;cH1>A
58;+S7J-9f3I-I[W0LPV44:<Vc@4Ff9dXU=9YX24_1:.dD2OQf\cF/5KH70g/1:>
(R^/AA^,_K(EO,^^0\)QSS)ME6O6A7N8I:UVb<2UR]S/?QMEgZ2)P24]dE=-2,?)
>+KW3UVb#7)AW5Ec(5+F@=MN__c:G6;0-gA(-Mbe]=84CCI[?IJ_BLAWc8cX(R-A
+-;-PLN<+d/D@L5Ac)=:IIW3L;C>]T_;DJ^TRV],OI-?31O&/3Gg]b?U<ER#bBRQ
c.F5:FVdUFI/=gc@X5AFBDb0Vd&_W7e#gTCM8RU[N15Z:/.7E^QN[f4?><Y;JK5+
#E?>I92IR,_TD>3RM=ZDX8Z]Y)V9PO/:OX3C0geN+6@?HRHUPScBIdTa.-f3<>IP
+L08=R?g#2DQD,-cc>(-TSCLS=PAW4SA_+N<-b7?7.3Le+f<7)/F2;7?(91RS3\a
)M8=3JgK14E9EfUN2?E(g7\18UAEaA261SdN?]>4,DR]4\&:Q51:VLFMGET3bdFA
J4=]N/1H;0&\[@#)<e7NQ_VeYUGQXNBJb63FT:OU#8=M[ac4\VR?V+cUM]0JV>fe
YA;8F[^F9-WdU--D+NI&,JM#7?c#.d9O6=6Z3S@5U6f&<;\E\aCGM?dbL=_FPg:(
82R+Rd/GQ-8QC1T?KLY[58:I8d=dDd:0c+>]P+JDTGaD,OMbBV3MgOV?55Z25OAJ
CH^YV8M,]&DR)b(_1Jd.A:K7Q:EGWIYJ/KR.(C^2-Y<f;46+JS03XYA3LL1^a1PS
BZ7-.CXP7#UKf=HS(Qeg<:GX#T:&N/E9&#MG/\Z\=VY).L_,EPdK@)(JSM6U)OF2
>MYY1gN&;/^,P\Ee<MW4)/b;Lf#f--V0P^^bF[H6EOE^8;T41\__YbI?=_C1O-cU
1.Q<TD03VZ&Mf&.^(5aDSLAZg\LL:2^\2K-VK1\AZN^.6@A73>,ICJ97JaQ>]1BR
0[=gf@DE,\4:FYQE\52e+/9<R_2A>DaIAZO6Fg0CNfP2#3<DR<T?^[X>(#^^V/:a
JH/P\L^;H0L3^M[@+>GAQQ1NRMTBW.].N;-Ec.DcZ3W-Uc-Fg,9da/Lc8GO4L6&S
gE+-6>V;8@+P7fRXdVZg.RCbBUND(RK1MFc.4E+/),Y__)2&8De.M/edT@0;U,<B
+ga9IAIB3Z6Nd+?U3W39PV/D-PZ=aIZSgXJeM^KQ/_B:<gfU[+TM?1K[RNF&&Ia2
M&FG?_ec3IZKQDP\R4PWg)MG\;Q7,Hg<.CX09cLD3Se7>?26^OC[6X^1B)4&<G;)
aC4XaNX-MD1S^dLOW<?J\cS]bKF)cE3aEPG#(^N\CGX?9&?QdVXN\&V>#@Ge7+R]
:7YVdZRb(/Q)EOQKf6UIaU/38Y[H#gc5b_HK&W7.-dDDB/2/PHY>9&aS;&8YXICF
PLadQ(Z2W+:4JBI=DV@J>>AHLdIX5Kd_4VER34M;C]f^:ESJ#8;6=IK/#I2GBCc:
V>_0[75>fW8]M+K\GPQ^_].V^[K:P@)?._?H.63W+0FXcG>=[ggW2)dYCc(@Rc&D
,1,K-.;Nb;_YQYO7a]DE4S8D?0LFO57((^,0[UHC;0^Q48FNY&fCeDafHJ;QE2N?
aTXRG)SW;YVg&gA38J8\2&Ff5N6#^^d.(UX#6:GVE;K6@2&Y+FRaQIM7,[S=e4@3
.W2dCCKN]])19+C-2AV9#^IR:@aN4.I(W9@R[(OOg4geUTbGCIQ+V?D&<.D9bc(c
[^#a0JRIA,a;C^F\;;PU9EO]9@LfdY63IOE;C7Jf)\c-P;_E;J#McIT]:T<#EgWa
3]Qg8D)BR,--QT1^DD5&S<dZ)<@Uc^4eFB5cf]I8H5-#L<6e&KW+?g5fH7g?0YUI
47TO0@L4G9,5U2R7JU<D>VTK5:7P66UL#6Y,H5b<,2&Q6YCaFWc9U5F3LgY8\A<W
\72:ZaUF-^9[B0dLXCB55gWS?/Q5cXVT/YKNgXBMRDcRL+H2bKU]_@6T,6OE0f\T
55J.0QYP9dZ3RWK?2dI.<^.5KgTC9?=8LL>2E_O_cCc.cc=3+2@VKP7W+WHU&\Ug
.7+U6)N,gC.2Sd#@=UcBTXdL?EY&6;)8V\-82PX,&DK+H.A\B\H#,b>MO<bF@8T?
)b9]JH_bWeVW895&\fO<EM65WY0c2.G_X)0A&((P72<f7>eNgZ=gXUED^,b?2::O
bFa24]8SXW@4L?aRH/_R+a,O/_/LG-LPCG^0bJ5d_]T]YaKZaXH3.@68>J=)UMc)
O#PgU=]aJ:?,I[@7d>@#a3\EBP=^T@<R\BTIRX>?4aGC9J4ZJ<@D]G<acP;FJ6>7
\b/T;>6=#=BXS/LdC]IU@24d@R.J<fC3VfOL@=CD-8_M_>=(eRbR^c-2N+FbM12d
3)e2OLJD_-&>,f2[CO0A_cCE??03?8#)-8dAY(9eS)7>3CD2ZL?FG=LBce>0d@S/
;CV-SdT+Z#7A?b=KQ5&V0CbdM86XKL_bN:9:WFaf1)P)8?gN5B0<7Td>,Ia,H@AP
I>#0/PAL\7PS;@9C(aVJbG./NE&4([KW&0X;11bEY9MO8F=1JY@FU7F7N&<Od5/X
RaR0dDQI[M_:SQCdaG@c]2P,PfKe(A+b[YUILOaO?@O+gVF0<]ZU/JZEC]42V138
^,AFOQX3HHC#K/XQ52@C^6^U\LWW9C0D^0_a<1?+e0=+B&P1YS3DFbFJ;d>VOa)/
L)>9LcMU1KObL6QO,7UYG4GWCJcV6cD7eR6QaQ\EQ-V64g-7<N&5_XdPMeD.XXR@
S,:8VW.L_G:21?>>-DOU^WTBU)Q_VYb]XBZV0I5eQ,/QKOODESD\5DY+f)YZ+@,[
E4SEN[YA<;=U5Z)EdWVE3ZMK#6L-Q2ZOMN>QdV?X\,/N(HV&_YLcH55,1KY^3OZ>
A]<&9dgg<7-8)C0=PCQOVTF7>IZ9ZIW5PMYC1>eVK1G4]-U8Wb^A2eA+T]/]ZEAN
-2^#AJJa^[2gUBXQ^@C-LKeT-WV+ad.<G^U_^LJ9]3=VR-BZO)DA3,cEEacFUe_N
7?c@M+ac=)CY,V)U)Z90:][<0AA:-YY+.BaC+@g\PfJ0,FXK+7gXbg7VBdU9XB.Q
?0BKM/P,VY+)J[f\01M75)X5F\ROcN0cdK3RWd0/;X2VdVf?VQPE8+E,/cBbd]/-
aFfVZ24@6gaWS?NB1+;Vf59N^UU?ZH7TRS<@a?1IT\fDUO=1E2V8\#O5g[0VdLC9
#YJ0N-+#=<Y96PCF6IW6/[H\R7@)\XS3?KY0]2LaMdb<:=>I&\1C#SA(\#\S<9J[
ITAQ2f8H,/#&DM3F-Od<fBcA[W/T3QN2;T//0H1MC:18.4-7c6Fa#&4#=+WeI;3_
S1MdbFb/fW@P,_(CbHDN2^L94,@2(J^B0G:IMONWBAGM7/\ZgX=38P3.,,W67Wf>
2B[]OgVLGM6PKQf>QHcF=SZ@g9gY.J#J16GdbP45#5Y7[I\5B13_.BBD?(3_Gg#A
g:[ZSf^)>L-)3V^N37.b0X8O:H@cZ3Xb]dbBNd])@]>S9XTQ[4=M)Fcf=5cC_KTa
^EE/9_[:T[<DL/AN3Z=fG>YRFG>?e\0.WX[4O4]3V:J?,VPH4T^4?6L05;4=DAYf
5]^_>HA:E?Ed7[f)4.8+PV]MX0LXZ17=R<NON7&C>Ze\1MCga354P?-FODCc8)0H
>?;TR?/OOE7N:JQTZ-ZJ/ECEL)K_e2+(GBF^WVS+^>3e]\RF>XO.DaD)SB@Y3B)7
0E1FA+7Ac/R-7\YT3U3=0VVKR.TZc8X:YKD0HL;R8E_e]TQ\BZMSFRF]S:N&(W@.
7Q0O,XM@VCJTVMMd?aKXH7U0E):dUXXO/E42=.a-1W<dGBC7=L-MS7R4E3_M80Hd
MT87NJeBgI:\B(9cPbH^TQY6B158FK<7V08\NH]0T)BMb=2&WU#d8118YD]R>R7f
9.cWd(,KMVH(XVd^X6DY^_Yf09;1+.^O4^#1eaJAMQ29Faf_e,UV;Icb9V3R_\_N
&U,R.IJ@<9e6d902X6VE]1[FV5\f,]L.[IC_EHZ=H.RWYEaVfZKLLf5fNH-RE16#
E#0[W9-H>Q)97-P6cOa=9:?<,3eGYP:-)&L1PFN[?fe)[IE^gWYH9WV5Q=fCF<[@
FZT:TF;.XG_2f_F3@74461..=dE9<c)@Sa@N4/6=GT-E>:2WVASF7@#Z1;@dSg5=
+U(WG1/-6PQW-7/#;.A#?aP;<O_J]9M&0;NW19#\A9:,a/c>T#X:4FVSRY3Y/4CI
c->64<#I&G3/67))ISI[1,T7f&If8VZbV3EZbV;@fDIGPFPeH@ePI^]Dc>4_?C5Y
Cd+842HW^3EB3-a\)dIZN_=g,6WUI2\g]/#MQUYdBAK7NgVbKU0:-CD@F\]T&a_a
8eIU/9e[UE#5S3ab=+DOTW1eYGTHD3(LgD0-E+:[bUDQX52/:?X1c1MWFeeH>T:W
I)\cb]X7XLa:W-&X9^[/P8(__2aC][12.9[Z8f]W#N4#+JRg<Eb#-EYf2XdPTL?/
/@G120CYdeW-131?daKCRb6B#M)=MD.K(8R[_0WDM?N9OPL4aYG&Y0a#TIHGBPCT
>Oa1,OC4F/C<cL02:P7^I;N=_:d=6=[6)1H<4LF7CIO&W?<=2#e3[4\DCX1fTF39
#XCY7,5JDX6RF5cG1G&3bTVAHN@T8DH3O4/@\=H?cZ=&PaV]4J282D>&XW6-P.\L
VBO7.E0&-W&LKWYWWXUC+^_,9JF3KfRWQ&3LMS:0WOdVdYN/\.afZfWJ_R[[b8Nb
#VH\CL&)OQ^/LCX38WZaOc:]J-;T]AeV6V;8^AWSBNG2Q<15\\dPN=XCKF1V1^;c
3S:3L&Yb0S0G&(VVP@H2:_KA51geM0H5;ZY?d6;1\T>#e,<J+Dg@.N),DV<=->R1
C96<)68Z4aaH)d:8d2IO(C@)3SK13-55@T=F@;eX(7PS=3<3HgFEE>D1bE>0+g\6
DF.[A&Ef,CB1:\_fVMS+LVV]X&L@82D0;;GGVG040O-&9c/W9TaV[&cFD,[6C[)a
:;NS\5P[>4>4@9JY7N?]bUWL.AHBQ9:A]d[25g=[T;(RI,GNG,f2-BF=EXBDed^/
dC?G<QQJ^39:P?TX:D@HP:4,SaKYI1]Z+7PNK<Qg&T+\QeB,.AEYUY1(]M()E]Ad
]O+:QIg<CQB=3:PYZ3X?T(;e-T,X<B&eR0D^V<(0b+If2R4RPUKaKIF6HS#_-eF9
D/JCZM:d4FeO2Q]VH7T9M[))(CZ,=b,1c-F>d2:g516/91ad/AWa^Cce9,L\G0@C
(;/&LR0RaGbIS<YE2WC,NJ,UFO34UgSa?DPE=DJ68U11YM<OCSW][N#MTMcUPb][
g+c6N-8(ISdDQ<JLMW<7#^P-CeTcO=T3>I=-E^K#GcI9.[baHJ^#MSV,^IDZ/[(7
TE=)&F9L3I2CO?fF6IP[RC7S<f8S3_VBbM7f36?g-X&>7MKEJ3N9]K/b4.3N6ROC
T@N]b[&[EA1F&B3>aUQ>b:_a+f<A2K.77,9L@ZP/_++=7PRX26+=-&.)WNF/QeR_
(&Y+N>5XRATUNO&E9KB?W741SSbC,AHJU9ZP7W[T(./=N<@Y82/5TagHW2-[DQHA
,dc[FX=aVT7U7c14/RQ\L76(\-<;^#1^.)(#_DRaE5,cJS/;0CRfBU)eTQ8O2VNG
d=)T/J_a2N/#)RZT^6KZW-W@&R?=F6Bc@ANa7(?.:gHb44Kc_>#J>ZgH9+L8=B<6
+<4KAFI.I3&4J5(RD\1ed^1Z2?#W>5-I^][,^9dXI6<RM=P>E,TC^#0J+[@J4acH
,3+=VMC-Y7\4c1\(/UZ?RAXG;3VYUbBAb,IX;8XF8]/LKI)T8PaA@;1-_(c:#MK-
-1D+/56LNJ?[RB8ZJ65-4A<W13N-g/RC7,YDgO]3c;D_=D)>Z:gNbNCFV@DdW(G:
Zb+@Se^d8WI2(E#DZ-=(1W_:Jf9W[&BG9(2)L>@<W<M8CNTg3b4fgHS(91L43>GA
YW\NPg[[Q>9HG7/CPA.O8GGC5&\Q(Qd?6.89LRU_>.<;g4W>KKV>P(e#C=#F2eI8
Rb^+e6cX+7g^]M&Q]&E&M@0+-]CdNGT+8:gD;3(:&eP,J3&U,#[;\O2V;UDaY[NG
b2G.:g(40?OHJ8NSV/Ra<K#J._dIR-<-LX9Ea9^[L=C>4#7eHRbMd=F(K]<0_;NZ
81Sf/]F))RR?&CUbaA2_N.ND>fa[/aKN_^f1P=0Fe^&5E1)\[F@g,=ZUO>.56W/B
X>JU5AZ+43:Y>,(=\=Nb],6X;eM?7M_Gb5D,&M9]6B^?1AY=e;9/OHU?V6A\U1P,
=&BT6E+DC)F]@52b&9EZ9MaV[dWMNRYWT6G0P#b9#V3&]DVA:ccdGMO+D5.AE,L9
MFQ_(/g^gEU6I,YN@67R2B26@:;Bgb?H0@f-9,EZ7M1<4L>:RcH)64@>b:2/]=B>
9T7Ba3,5aUVc?9.gBVc3I.8_=MKA<=faDd?M;gagCZQMH^V,cGc-7KT>I41H#KK6
aG19\]Fa5E8M3(b<,CbXWf;g(U:P0?IDL=4fJ+6AL[VT?UGGVI)3&ALP39gF[4RA
V>=5_-:Y@4S57Z<U4ee^F_3?LLKBU:QV>(C6L8S>O2Z.:6CA[5@28(ZE9QF,61Q3
Dd^B>/\c(Ka<ZS^^C\+770:6;PM_b)Q+^/Je\N(bXKea0_@@5+:>e0c@Z6cFb&b#
ag].K<\XCg3_J[AD:=X60VQ)9N2KUIN4N3bS1[(TI,c?@+OMD?ed<O:\))e^WA@b
<+-g)e4=XbdSD2CG/,#SGY<<><Q]8>ZB;,^gVg2f+IT2B3H)2G5BX\F7G1DOf+X]
b8dfKFBO,WHUEfCE/W=3^01cY:5+cHFK2FJ2605]=DCJ-.]7V4Q>E;7d=51Y7WKP
]ZN>YD&/=^,d6P_2XETg&T_?SF1b2C1;cab,>Dc3W,+AaHed_Ne7Z<1a+^cIKI29
\0L]M0;38G/OWJSd_a>K8aS)IK5:Fc?(Z;<EBL8XW-e.D-,Td]Q0W@AEY_]b(3E1
T=3,O7bU6YG:G9SQS=^C@cW^8C@Sa7V7\&N@H;LHMT(TIZ.TE9R:R#R7a[MUDVa+
4R+dP[3<c6FWJI)Ce+U5cQBgcV=YS38,A7eRaA[9493G#N:[E=<;^I\f@M:a&4>]
-/9)S?OHJe9DPTf&HDEfF87=^UFM+7fQ6cb0V&=CaCEYO(5bIA(WU(5-(RGJ2gW]
UQSV,2.NeA4RC=g-HXc-JIFcG[Q,)e&FVI:RA-R5eO5=MS5_^f^fKZ3+H3/-ZaQ^
^=58R,)JdU.ZR+ZX=O,[b=K4,_(aB)>S,E(J8WQ-c]abERR7#\5)Q5N?VM4V,T8S
8a+;Y6_;YY&J)OQK8ZRKC4\eaUO;#fbEGU&LgFBfXR[5c]MH[V:X[.VV[,UIEPUa
cb(Q95Q/4=b<c,[BG5Z,B.\DYP/L2B8H@[C93;O#JWb#KJ_>]./b^^e.2_(6S-.H
,NNSd2.RE+:JO660G6:#0b(ag6Q=)aHf8#fb55HF,JL0TfO+0B7OX3g^A98T(<37
E(1L4XZ[2>/1=d_4#9<FbPWZN<136;JJcX2IEAT_1&fH\[GT+X\^53.IITQVC7dW
83c9Z]Sg6Tc0+ca[7[/;#\\LU9/;4YR2)>AM/J=4J884:^;R3RG1&WOgC0HgAg47
B,MX\N&b:L7&A_XN72&ZET6Je^^CUU^1-)2.7PMLW-eV1IR[T.9_Ie+.NgJeAYGI
R33dBE6:eRN?G83D4PTI,EHOfWJd6UV3<._7-eY0+@(32WS=PO0RMB\ZZeAQ.\(D
EID_b\gZT\,E_<>:6(U(LE31?H/-P?L#;=?JH4&^Q8P5]OUH]9YD.f\P)XLcbdVE
\^a_98)bRCN^=VTVU^BRY]7?0RC1SYEBA+9?R>g]HAQ8<#GI<-^36;WZ&(E@53\,
dA6+V-ILf^]JN0D(/[:&\f4_:5/3.8TRFY^DW:M>I#a)V2aUf^KBHad[0fH,)O6c
IG3:G9C)#?W/FE/\#GED5b#DDRSFa;AYeG+@g0+PdcSbI_[LWb(f)/3Pc;_C?e1,
,IJZ>G(,0IG;FB/K<,<7)@a[=fTP2]):N_<AXRL1?CRVR3W[CW9BXD&L4=O>Z<6\
EB#2Sd6WSJ[6AQSaLK:P>F^UU>LUVC1[;<8E8d<I1TCd[Z-BYDJ._gf&J3BW3-L3
L9ga+_9Q+=TNP/,7JLce9>bXHO0-\@N#9_G7A([U>/@2+IR1=8RBSaXDE@NL#;L=
;#P=TP><KV3Ke;]#ebcUbMF=V>6C:37&-^SFS2,L)&KXU.CQC;?D;ZU824eD>M.-
2a;-aP7]B#0F#b:7ZN2bS:Zb30Kc@Sf9>OFf-/@@Q7L5C=@8]89bTEAI7&-_=<Z<
FI3L(+6R-66J,JV+L7Z6RCR2g+6+A+ALNG74]e#7XO7#N7W?bWNe?LWLdNVGS=T@
_ZgC180a:eZ,.(eT>FZ^3<3@2MaPH?>O.V;11;<8a]YI=7f^B?+1RMHTV.f.9_&+
9DbE[H.bYa9O7g_IPEK]-BR.POY]F3.[X8DWdaWgVN5a[^2U9A=]H:eVeB2aaGD0
]MQ4J@4B,@#eU\aDaUH2cL;,=Z4/Z8aB4.PHWG1)Q:U8-S?Z0UVBQW=1eP\bFc9L
f98d&6(O=-AVH;M/D<EeF_D]\]fL\cFLL]O=,BW3MY^^;Ife0LV>I9[+6D2(X9<4
)Fg/Qd+e@LCV/LF=TI331LQRKIYG)G/=UgLG6Dc1\LI=NV+]fX>0e[UOD^)119SB
3gaF(L?BFd)dSHVLdR9U-T8<0_6dMRH\f=H=U=@K^],\8,#c4F+,IbB6/0]#6/=7
79IHZ9B/6]T9>NSN/BA5O/d8YOg/F3egNZ(f7,EZ2^)HNN1=EMW/^;SYP2Z)bHc_
C_BM78LWSgfVdEJTBZ@fG^J7)f4=)EJc,dH[NERHGV=UZ3_Q@3MX1aQc0e10S2SW
&0ZgKRQ>Z#B9B>9LT3dO\U.:[+[CV\K_3CV65_YB9T,X&\-5eVc?TC(2R?1M3Ta?
0)?O4^X745/ONTYE9<ST,f1KW.<[&03Zc6Rf^c.#602,Q/(+e50gf[(5]OO&P?+5
9<ZePK>G[Q);))1Y<92(O?fD;U#0]df]M,,5YLa@N_D3:N35dKFf#J2J(5)XaG/&
RgJAV2DH9U5Nf9NWa?C7MR>HBCT497<T6&=9f_A<)V2<2/F<D/]RHSAgJe[PX(\3
fW\52EJ)[D5fY].d:@C91+2+AN79L9V>B)5:ZK@\S,XBQ^+aW5Y^gg-;Z.V,Yeb[
+./)7U6dJc>:A<.VG&.V#OWd_[7GEVM0B_401aGR..@@ID6V5@@4A#dIXf2S=>9g
O\[d&+A(>QDY+VQ9@,g<dXEAfa)XC>CZXfNT9YX7X[<Cc=SQMJXJE/<.#f&?@WgX
;3IV32QU\4<CW^^:acO0,EVZ(_Y2#E6P;LI(bACeA1=O&e5Oba:E:;[a)6)T2FV(
,<I^c4UUERVG.Fa>E96;T/2gBLEB;V_.K8ce/GDaM<&Fg3:I3CbgDE=6=)QNUMd_
>@d_ED6,E1ZEUFKZ24CR:=)(CQV^=+#.1]L:X\)EW@?X_AA.JVfX>H@)Mf&]a)J-
=9HBT&41P-TAV+5EIX:a&:?/,g>F>.P,5]XAZ2)cedCS.5KL&;JE+TC]g>8BF;A.
-/XJ/>^H<@KPa^A>+UdH/\)]:<^0D(R[C-@N52Gc^FQ+Bc1<OgD61B5(^b=UU3W^
3>3+Fe?f6S7CdL&DVdW/D9]-1=D?S@U1cOE>C+?@[RH\X>(/8CUQgU@ZN;cX?93T
f08FN^JKN&XNPRJS9))PK2+H28=M;e@:W\5HP-O(H^B)\ZL&BU=<9,-<S>&C:6V4
YRU&59NAKL:@f>QNI2>L52C/7b)XTHK(+&SB7H=g+LUMe,@<[U,&][W1c]?DAW_3
#B=EDMMKRTX7KW@b,dJN[-ZMGXX[<7B;LSC?I3+:3]V;IHYeL@BZ(BA(H,:2]a4L
;I@@&SCLX#-\3=G&62A/BBIRQD\\deS>3_53V(F,VTL?EBY2cJH3EeaAY(Z.QWUY
d7J/D&Ma6D@6[dA3&e4BZ\JP?PY<4AKa4(Z-eNf,W54&5cNN,J5P<Ye9V9gO_5A=
4(3XVea+MXU?\TZ>MY^^4W[ACS4SP,8OD-:TB<9;-73\;A6.:297SLO99IQ(6a/7
=2.@X<geUfN<09I\2#6)QQF[_)<EGG77Z8RCK#G:PF;4(O0FbFL359@S)XW;=HC&
])RJfD4TW(SC;S=?F__/VZ._8B3Ua)ZN:GM;b>:W,F2K573?,@XT11MB5K^\Ae=9
LV1]>3+1<RN[Oc2-JS)eZK(cf7d&4[f?Ig:b?a:1GXLD^>X2J_KW+ZY5V1TZ0]4@
:RVGA-X9,bV@3\BF=g-dR;aJSW6NIQ#JWK[f5Mg[-><DU;U]MXXF;Jg=aUYE[&7&
_\b8]PI.aPb[55#EaT33YJQ[GV;9,[BZ63#IY]THWFH&SL>-3]9#)DV2.OJ(NaMD
J,Pff&0>056@)J_0L_GZMg6(3R@C=0B+LTaT],I/^CH/XFALL(C\,cNcP\O8R#78
\ZU,&Q3?XL^?SLd5a>.g5(+5,cG(dCHJFc6QaA3=S-^bH9;W87g_/IZWK,-S?AH]
.\1PHD/&O:WVe_=:C@gd&BH64>>EBVQ\;+ef(U+JgGX0Tg4;DZ,:;A9Oe4#-;F^f
O@ITQVJ;d]]fQ4=2a1]g\ELZX75_T]3Ob8](:QU_&K#.I_O\0RUd@):5^#5)<94B
45]ELAaG,7gLG&7Z@DSUWfQa]ZN8Y>GMbRBOHgO>_e?4eCISf,aGL<H^@WT>F+M6
GT4)TP@J(GN06G1:L2@H2E6W7S=)/-;[UAV>N??&8MUW3G<AU0E,fe9Qf=,N9+DR
\KR+OH&5Y81c#_Z<@9R;]OCFaeYH)K=+<;e<&+O3<>K9c)U\aX1_PDQPaFM9/1:&
J?#J1B#_^03R&DYZPVR+V\.69@GD2++SW-3,.>GHZTR@.9dCY\8QU)LY#KbC^.=Y
2dYEN<)50D?J6FYP+GK\XXQS&1dT4eN(9+FMY\52bfU)CX;K^]1YdO)L0(]PCW)/
Ag7K>b3N@(eOC3AG>fg.]F@.6_KVS;#22I</56cNH/M[6,FARePG[PFN)G2UN(&+
5P/K4O/?O1;d9\A\J0-M^)K4cMMKO0K.)MS+,gd:?9X8SA2A_WdSdgcIYTec5MHI
=]ER8Y2BKRLKH;_.4)3]-G)80//D4:gG,fTCdCfGRKDNF(DGaT++R(A<0OMGJR@Y
MQ+OYLgFF;,D^&DE?FN&G>-,7L@+8IYK3]I\D:O2feG,ffg;QLcb/@B8ZT[^EPSI
.:PX:(cP1H>T\c6=BSS&-9F9>3(WaUAQ?Ie^ZLU>1K29CFLd7DbJ&)PX_UFZ(SR5
4252Bfd35EI2B+bO9.72g+<P>]CWB+b6A6^EIM^SaBMFg]XLe0?a[_(:1.d1G+TJ
IFI3b0_OM/X4aTS6G]0IEJA4I_1Xd7&KgG#c,KAE.5+LQV>@EH3.aQE&AbJ:)b8M
f2CTE<DTU:W7.Qc.+N2AA^JCSIbUd9?\JYU?0a^N\<2La8g[^56UHL#?W/]HHaRI
8KTLKGUJ2H4F2M;X4DA^^dCg25@b2F)K@-=5fP2@[Je#._Qf<+TXARc\>FXVX2)3
VJE4SU<(4@^#?cGcA8Ygc7AXOUQM_U=:aSYc62MN\aQ,]eIKI=1OJ29Oe)M8-G68
gRJD?V,SG,:U&H&aV-Ye.c_4.UQ[^CX<3@H)f_O+;]9.R7XX:X+@](c;gXT6::VV
C<X<OFV6b)dH_d#08/?eJPWL,:PE6?J;\B+RGYJRU[[8QD@+(/N>K,03\MJ<5g&c
f8];?;,F52NPQZ;Y^J/4(GTfU/eY)HSE;Z?<E<91.LcY57df6[B6B\B,EQ#[.(2G
\V:^H9,3=G#0F;X&JXV;778DbT-U?E(C,3KL<K0J7RfANSQ6U.KfQ)G0TEg_]O9a
\\60d4Ngg=Ac,7ORZWdU11/+^>V1a]GbYg)dX7Qg/O8S\DYV@?e_VA^8@):M5^48
<6HR5R4eJWL,(:6^W).&]E^.M;J5_?B59])]RU?P?@BI:<W2fA<5a^APEa7A(\7+
b7[5X04UH;=G[c51cf/.b4]P1<-[+[JS=.^e><.J<bT-P,I@T+1\NXTQ&aT5V-e+
JU4]ddD-S.3[WR#g^QZGX.4Ga7RUc<V/;&d9UBaH05:QE@R,(B.>dOL=(dEX9[E[
g@)d3?S.Ja4<_NZMc-]f?P^V7;SBA(bTG^JVH&0TS6&M[B;6Sa3;QBCbXccDDbBH
<Of:DAZ)aDW6E,-R,TK]I^M0Y34-UCcLGIJY6YY2Q\28\UQId>ZY@HGK3Zg@d7ST
?)d2TQ\2[LXTU.G,HU0Le/NTNTR&+V\CARZGW#-Af7-.-Xg^KO9O&:#fYL-[7^-N
:?&g4dTK?BX1P8H5)0NL8XY>YNQAB>S8#L/TNQ/OWM9\B#V4(37FI+N:K1HF0=(\
e6,)G)9?]=d^cQ<Dg-)<P5Na6+++8f0Ag-\Y]_M?N]I&3R@:(8@0#12U(SKbgSEH
@KR_G<fYO?=\HG\->@P4ZX]QPC<XS#8C3Q?(fgOgP[9&I#@L]MNIV?=SB\PS#^X/
7J2C-2[-4+cH4Q\4I_WL.fH>T3BO73?3&-IOLZM=d>afeI^XGf\?QPN;-9cHM,<J
4)E;:7G^J;;K3VH51H[(GKU@D,C,._2RL&&/aXX9gXUD?H6g5.F[/Y_7_O_-GaA3
\Md@13)TS;7JV&5U8-WK4,fM,S7&gP>U457a5)HPFI^7W]SVQ7P^fI5BdU+\eQHc
#45<&&ad>3O4_.]M&=T]aQAf6T\fN]S;\XV(2M)HV&OLXM.4(aT2GSQ9(M/_KU5I
WPJHcDD[HFA@2JQ7>],TaHI^dZ1^RFK>8LI.G5agB^NR<V3B<DV\FBVDHCNcgbV/
@_,8XS<^W&#bU9V72Qc\6L:OY-Ff5P1H-=B:Scd/@B91Tb3&1.[D]5WSa5dC94&O
U59:[=[Ed,[?[@6R.;F:28;4)Of=4J^O5=,)ZWZ.Y3>VWV8Q3,a;>g+5OdY--HDM
?D:W(WA[:,<0;>GTNC4(S)56bPaW5.LFA]-FFFPJ?:#E9Z3fH0RFb:cT>V:?53-=
;1D<1g4X#ABb?UUZ<U&-1@PSbfIXbX<HG7Rg+7B8NY]<,E)c>?@XaR)&O+2]B9,[
_Gf9#=[A:b+E704IgG6e)W_d/Oe1(&@Gc?Y\1^eF_\KZcVI#]E_8bBO#)4-)8C\:
_ZR[fP.V_@KVgR_0aR62ada?[Q^_0_Zd_@BE,Ie:a2::6g1M98E_NS<>;NP5_@Jd
#X@(X(BKTfF<Je#Z.=][E?^1RF)aQ</LXGBJB+@9C_7RDeV.:HB:8KCDANHNc8P>
^SBPUc)Xbd?[Ld@/f-Y.#X7g9U\OU@;bW:6,61)?c10d8Z5^F]LI3aN0Z+S&K)_[
>FJBJC]3bU:8X.WU^NT1CC7f?.>X&X,Q3R;eX6A\EQP/)0J<g.6/61S8a@#:YBc#
=TcU(:&#JR9>1[+6FT=#QBV0\62.WDOYZg<50OUR;YD[N\RA<&J1aDg175-)ZOWX
)9eE2BB2FGFEGOCb?4X4Z1#FC5.,5S3J<PA2d@53@YW(G?3=9[W#GWL?f7g0J,5V
=>3C_HCKOgLEMd3\_#161bGPF[>4M?RN/Q,RI1/1E:JG#R]NB>+]Y7agHW@[G-K_
F+9DP3=Ze-RLf8].L89R<\R,C1e-@[Y(P\6UD9.A@IbYW9IeDY[ED/M5QM^\72)/
C8.<>[F:NXf0F\]?a8TYVV9?Y0_d:gc[#[;@XV#(_.(4F8H07@aR]QYX.FSVFM#O
W2Z6R1S&1O[;caO0>bZKPcX(ZS\(_b\^IQYM1UB84cC)@IA]_ZY:_f=F_^-d5RgB
PD>[MU-NM.2.6Q(UFgJ4)ZFX&=S2CKXeRJ>?U?P=PMc#+;DB&AU4C]g7eP3Q=^Lc
_Eg^>4>aIf<?NX\[)MYJ)OVIEcc-Xf?KTNC:SOMDN?EUT_DXO/cP3[B@S/b]M8XT
fb4_8_>V3Q_f4:_,&8=;8:O?[39cU@M>GNVQ4)bE3C-7S@c(M4]4.3bSP)-@f8+,
?FX,Pe>1dDXfc&;HI];_aUgcW)8Pa-LaS1:7F/\dWF2f=cJL\H4X[ZgH7W.A4K5F
,gC=MI1:KT-UVH?QC,5YdOY-a_C\UgSd=T>YOE(V_8SLQ[.O0)X7g/O=P[WOINXX
VgVOdC2T31?NSX[9QYb51e/Q]?3)A.M-N#-e@3@5@6/dfY3LH?T<X@aF=9LJEfI8
^?4SPaBeY-F[];POXdSFLEH-UWTQd<4VJ.(FM?JPE3J8B1S,Af94BE\E_Wb.Se\,
JQ9ZRA4Xg2RL.V;J]J]0QA1L:8(7@Z<9c)?:E?J,GXFPKO104bPaeL0>ESf[=BG#
_^MG-L0/7)#+8C(N:).eRNbc6gMV?3SBF7Y,S0c>W1E-V+]#PKN.?B)Y=g8Mg[(C
@\,&QfJ)g/F0^&aYQ_T9NH33IbOFLC&<.9156-(ZO?IC^P6=YY,JeI(/G3VQg,>&
5[4e/1671EW1/3e[)N(gC-8Eb>Y@=CX;@9QIS)HCe2gN]ZKJ0#<T#I-9/P[+4IMH
)eF[g^H5C:REQ.+3CGP;G9(K54?7P?O>DZ?D&0(V9UNY+983/MKU>K2e4Z.85ZW?
D8Y355&7a,HJ&>C+W6>\Q.#GI;APRZIa;Q>]5&)Tc4?65?B9Vd]a9+S4EVQEVe4&
FPEg3P+H)HV-e(QJJ?JfP-)gbF81.fQ=M3-&=I3HJ;#16(RZ8D:A/>]#SZ?#D;A(
/FYO?XRQ#I<6RZ0E1FMV.Y27/S:PX>)RG5aaH&H;IX-O;^H,\^[7Pf4#U.DZVE,>
b^+AbX),K>8,EX5<<:N#3FW)PZHP=ObEG\@NY]HA2(23.da4dN\L);#dJZ++5eaJ
>AXW;W-Y7F+<^g\TJ5FPRL9IdC05EL\UM_Uc,O[d=H(U1d52DSQO;6(_[\_B-3-(
b&\@/2If#+S#.WW6#1^bN8#M31N(cI:FIEE17R#W\L^VN8D<a15Z>4.#SgH-?V4?
e4B/Ia]&d8:(OHYFC;?NKG98O@:1C/[T+6TRR\929]O]QS>B]@[N?JfV@K,:)0,B
&.@KcdAg+K[_DX02Q7&ZYR9e0:_,]c.)H,;5dfHS\GS.ED#.J8/3O?G0[(<ZdWF\
XfXb.((@@M#YV9]0@/_0=/@[,5^TJ#6ZC>,R]faZ:EBH(V(8fZLWbbd]Y2KH-ATe
Z/bMCMFGK1I>_cg&6-0e1]8F.F1NHC2QMV(a9.J,f^ZF^XCE8bON+/9E>1EaPQW2
cR8FGOR]f/2?-cg2S.]^8:_VZ.e&S;;FQA^NCb7+ZcER/4AK1O).7PGU5MB-(\UK
CaIB<+@.5+X=K/E]SA5=?GFOUg^SF,X<P7J4-TH,N8E]FV&HJWD(5I3[^&\<Y::O
YdT^U.9W-0EN)_DPDcE_LN>T]Od^2@T2__S=;4AeR:O47GXB[PXG^>[3WP2O?dGc
1&/4X=QPVg2?_:I[;?@cWX9@ZG);=>N)(5/fcIB,gS81?;_N.Y.45?/I6;<5eBTS
=S(Z@9(^HgP3De816:RCN?R?&6&CbPBL5W5S/eaZFC09<(8H95BMOb>RKXBGVZ6&
SU2OU&18>^_FRdK.HKeY#Q.:HGVMP2SI+TRd^6?Bb6]82IaL>DG_&LB/6O;gT_D(
#RO6PfFf-<EEAMA99>BHM6fYVa+S[UWQ6^FABbcbAdHTUb.I3K6<5C1+/aAL[2#a
4=S4#9eI@c>7VEJ4B79Q@+P^dc,FTTA7Dd:<RK1Y>,8\-E2PO:]PS=E;Kg@SgE3K
A(PDeQEC430J0WZ2#b?^.UG/dW@e;e1JY#;<18]Y)Q(fW@MV10=g&[6KVK1@7Db<
5&),Z&T3A-a=-;aWPH;5^S\7M..\bU<PI7Zb2D2e&OSLRDMZ7XK_UV?-5,/=EA&2
I+eC>70YN_NcCG7;89\V]KcTA\A&4/dg;TUWUK0CK&A)dI+<5>WI-gOb)5K&MNEe
1KTA@L7[EP1ER/C=3W@0]cG0@F.=VKTF9edV_H_8V?UKAXL5A901W@#VQ#([6]VL
6:C=IXBV7:QPaI6]_bS4Q1d^WR6,HP\S@F+1gA_eA9C8A3C<H,&E=3.#-g886fC,
Z9@94&1c>^Y-C-3,@f&<.7VZE&a=1N:3]f/C4RS@24[:-I/>e0<?0D/D4;(;gVLg
4#FU/<MW]Q/PJAgaV))JXC;BZ<^J8IV1G#=#R,f.Q7RC\[?fY:[g->Q0()MZ(;\9
1#2ZfDa)O>&IU2;,a(VMR:e0c(6_7X0>.eWMgF3ONK3.33:9VM[B?WHAZ-8c6^?W
8X9HTNE>0F/M5B+EF_57MeZ9XWH(+WU\0J?=f/+[UBSPV_CIEC#/?d?TKgQ-c5WL
d\KM#HbT;INGe]c256UWI?SBRc6MLS.bV^L1-H\T1)@PPTUCH:_WRDV_AYRFR6F[
H&]=+M3Z7]a8bHf.1DE8S/E,a/JL1^BFE_1DY_4,^&QECJ,E&ZCE<)>ECEfH>\a#
[,1DHV/P(F:1SFD1JR=f/T6_1;5V(:B>fNI5Y[KL)JR4+#F-FY?9F3#L^1)K_XED
M&a+Y4PINJ_M-I5U16=UU6LIVCbUD=(Y]4aC_<5dCA<[T.Pg94Q#W.):7g94?BVP
ZZ+^ZT7FS#fR62(DN20RWNO)/M3(9<QZL5Nb+4ULRQPJ1c=<G5N9;c^b1K-9TE0E
OKc0#J;G(-]2RWb]GN-69CO;<@IB;,\AS8?d3;1<6;Y7TXWJJ,61S+^Ub;e-5C.a
9ZAS(CJbIUI;5dPCL[.2SL)M2[2f-4b(E:VGD?(CI6S[X4SNb17Y.Wa)c[dS;-=^
(#@gCLBQTf92dT/4cY,(I6,H5A7BgS((B.I_+>8.E__7SL=<+.>,R=)V.@8>,^^K
O](G,2GCL^QMB4Ue9^JfL24AGI-d9LaWZVQ8,X.fYPKRFX5BTa)==+S-A[EIMdQf
fC9&&aV+RXR68K]X3-[KVC@,T9PFA7\L0O:L,g@:-TZaK)^#T=MPWVVc_VY#?AD+
>7P=_aNARBDeX6D70RR4a,C(17NASW-<QfNK&RQEdK)<&HeFZQacFd_X8FEf-_/X
E>b7_R6].Q(E[PV(>QVG_5LW&F0&,8P@VJPE7gTg0PFV-AL9;;=#PHN&O3dBg;V3
7)-K0aHEHS_DKf:gT2_E,M;KDC.]@B-d3bMPRB^)A)@>F5F+>DI2PN17^3F1AT/W
FWRD;0]GNX:0,dXX#1D55H<T+S=(13OId=<6aT82]P]23aHT^T^BZXGOA1\OE.H[
A^S-g.0N<)^9&,5\,EXY^gNHT<YX>a0>OFW66O,/M#e^SVcgY;E1UA@f,-HK7[+E
I,>^V,C5<LcY(UP&RGS8TW@/GMcO(bUZc+\Je=R\G5-EBHbVP\/)\)P#PD:A-bJb
6IdZNZ:1T>>GCfAM)3Kd9;REg+O+f7:PH&NEd<3U#P]T^,<(]3X/_R(T\0C0^@1#
cX@/7P/(JgVN#];>=:ENEY&0<:9Y+d<E^-a;5R6DVJ]+?PP]B/dC3d2bARS0RT>N
N.F)NA^I_CUF(MP_6O^3OXgMbHIXFD>SD;;Q^Jb-GVX5^Z4fc\S=;_L?X2^,#L&T
;JfDTVeZ?d:Da[IIPNQP2^\Z(=YH)3g#E?J>>9dCIIf)aIZ4FELCdW7/&<Ve[5Hf
7&(Aa^_geQXcdUL\_P6IK-6g(OKR@5-0Hab.dLM@Q-<,40F<V581&A-<TYZB^Re@
7729bE6_5Tf8TfO5,Z<GJ1J(RB\(Z;ZEHJ)30+&[DUN1L7SJ7_>0g\?@/AL))H;)
6;SgXfLQ1@8T=//PYg[Mb^e=;Nc<YZR:CT,_::W6e>.+O.U#DE27FW_P2\,aadJ#
UF.2IT1D2.(GE-YH1Z2(Pa]>81.KcEbKTP\DAC[RebU?I#:S8BfJ;SK?V[X/SR]=
FH0M+[=U--W?/,]Fa617YdCQ7BY0AY:YWE<AAJ^gGLc8A5_edQ]CNX/I^9V8+WQ#
D;N@P3d>d54gBO:8\IYKJ:_14#[eb_\Ie445W)eT91OR9SbT>(.1@CQXaOOU93YG
f5g#U#<A&?O>7UK>#3O-06RcG0],JBVDTcLJ6BW&1ZZ[^QD[G[-2:Z?N-LA?FSCU
7.c3a4D[[YU8@F:AIL2E:4AId?\&&=R)\473#K3[KM2U5a9D=&FB(^TE2H#D>)8R
D2&=TA3KWCd&F_)gaZUIa/<M+<Q5,2RgJ@=/Dd=FaYML2f-@7U4.VKW@SFYRVV@C
IL\>0HW(?A/aedAYXe\cg?Z.Q[A-b,PTYW<[7/F:YS_USTb6FdN>)8_T1N[g2P0B
P:E.B5bG+bXO27>L[15A[d/5R_7CFQ#3_#5\Vc^@X:_=]be9\U;=7O_5M1PH)?e8
Ld#VF[IZ+_GTb2Lb+?5cK.CYG?;+JX6gWCE_+/X4T3BFD7MGT(.UH(g3a9RI8&Rb
LL(0,#UJcP\;c4[#e-5;[LQIDD(_.SQ\/[(.):D2X,.R2@H^W_eDMb2),X6^0R3b
/e/59eUU+B.C4?+;f@9>)W5YY:),I=fKC_&/3dBOa[SVPXPSE8(c8WZNZ=00^\_Y
7UKM&]]BZI[SIA(=-J^P[MG3[I^2D9B=9V2BKU1<:/<1gIR^2N;UM1K/Q)BWf+HW
<1KCMN57TgGKZ9D?O+4g[:OM&1(f9M1^];F,,U,A0eC2[\(ccH@6EW_<#9K0HYS:
BO-[#KAX]79=(ZJ;<&c6=]aa6/0cRQ6)7d-SR,5=12S_G4IWZJ&SVVb@2a#cRAZ4
+5)G)8><N+8&H9M^<fG;XXX]\6@@Q?[/FAe>egWW>EOK<-4BGYP--=CI_c3L67>4
FLA&)PUHFCRY-8MCA=LCVdNcRROTPOIZCP)43&75,_++-76X4D3L.f86N^]4N\,A
0SF5W@._IRIea61O+fT:XA.c[D;WD((bXA=M)K998R<R)R<gB2@CI5)FF\U,J(:5
/_H/#?8ea^Sc6<SZY<Ug4)C^EJM)OMSQ23.XQ@\W:Ua6.XRKfS2V\)7eR_>;d&e7
7C:Be;a+3^E8X48)_R,8,HI9;5X,g;/)d3=FRgaD=Cd;K)2;0GC?3dd]NR/8V/5W
Z_A<M<XCdSF9AS-G[4E#LM;edQN71Y_S=gdEZcd[=.Kb;HJMLCY:.bD(IFcM56a4
,gWK4N/S]_W;7R/MYg@90AVP02AK#>O^.A]^PM6UQOW2\KV6IHOD=H>3#L0>gMYD
^AP55&>:)_MLZKbOgTC3L:VfBU\_G_N1L_f3;Z9?-&.7C,:_?eTO,8#CRJSYNd+1
@^d<1b4DL5X6(/S0W0CX#1K124.5?fJLPg,HD/?6=S5&?\@9f7CJ0L5IGd2-K/4V
/OT1T&KJZ/+9<3[DFIOO(#Z[MWK0Q>O14O-JX=]FgHbdQJM^.K]#(>M;(JgRGaY)
cH(g6:MA98^,f&#N,5W1DYY_b]S8=\9T<a84a2WEMcG,@&6K+9Q\Q.28Lf1=SLNa
5S)T98.]5F-L_[]1VD8/#D?&0Iga>E.4)U+^QZc<S;R<WL@DE1e@[gW99C59b7D#
,&-EfEK21+<)?ROQb]SDPN0KeaDYaZ=?N.:;#R^@..-,<@>#9@MeOJC<>SaNR4R[
a/VAC,#fJQ^UIQ;#I9e04de.+R2S.9aOQ>5eD0HId6=W</]RVUSH;Ed)\f:E.-@Q
Jd9fP@-V+\MOV[bY40VP(VfDI>F;/_QX>Gg:KaQ+cK/(OMUcb/LB)UI#dEgDR7LN
Z+E1_DAW]?XRDE]\Qf[U]VdI/?;H\=I^&d\?F(eaD8eN69Ya_3?C,P5]W)+8^NI^
4#fS,\O5aEc.91<Z4)+a?dB+S+#TeLLLf\+XH^B4f:21//#GICbb4/fB(Sg@>]CV
)PL+G9/(d;W\H\WcdO//;MB#M6[\<^NKGC;^F)JJOgZ.H_6^TF>_NZXIJ:0.ZQPX
S(]d0fE4LQSEXRE>3R(be;)S+\eN>DXC_;(dML+:a5=bH2@E(3K/J?-K+&GXV9(T
7cc3>B7,g(&[gY]:f-81c^+K>DTMH-;^[Q_0[SPR=gILbCB8O(?06=gRT:PRZQM-
W4KR)Z,^X&^]?YCAVffO6_;C9&E--(\[LZ#3P&D@f\_b#]eacO0K8LKS63S&Vfd/
WU@NMPM94-^f<(F@IIe1[1YLJ6#U8&7=LV^RF)MBZRg;W.W:EWK)+4S?Y0Kg3\f_
=VWHXVWULE[T3N]F&72HaC56X.)f4M/OT[[UV;d1+)NbUEMcg5B2YV9KK[C9=^ZT
QZ@R;Q>8?g&D2Z.9M?Z0F=;&DKCa(:._@>B3,P1f[NB4)J95?Ga3?;fL-4Oe3bGD
gEH+5:3bQSFc6I?NFMa=-]0KaD(+05eB[N0BRQ@>Aac>F[<Mg/_g[GeUSec42_Y]
c&;EO0aZ6Y/fKLN)]72&_900Y685-If)f],9_YYC-S+:[g0-X9<7CMf&@^bd=1a\
Md83O\\/+FNcbD22(_3VdNN#0cN[9+^O^&7^O4?N.5SbBZ8:=>1X@Ma;C^#K#)Se
B3,\Vg(M)+=2BdO3GX=ZQ)a/X^<eCdT1c,_D_>Q1[]E.F>?65Sg(X:5.,9^RACe>
RQ)(0;BQ)-VBAV#L;Z[B7HdKH#W1<dN]?8^RRV^2CI>>g5OA,P(7?O@EdZEVCYNX
1QGSKaeX5<eB2)#K3.C_OSVEDe_#@EcKA(c+J2F^9A2\_<S+B,R,5S;5R-[S43bJ
LAgR0/@O5HUE+AH>(8PbgZY-EI6Y(=.XJ?QbD+)fW06:3&&&4CJQF/X2ULaP/V7W
gP:cU>Z.V_RY?fa0JD7+,.CBGY@C#08>W,Wdg4;UZ469KN6HW6G&Z-PC)^7_Wa),
UD\,ZERdC.S7;ePWfa7EQ6--bLS@1GCDDWDd0ZH_-J9U0c?bNe10Z2TM>.8W>=/I
S)@9bU8LG0JRJT:aJN(Y+VKA.)a,5?1Z9Z=_NS>RMZfGDa_XM/e0E-#+A7/d4CQY
^;7a[FdXRFK64M^WW[T\A3>Y4/BbE[0M3(AY6.?1cI2bFW=Af#;dC;H8.D;0&6AM
Rg&;SDZ.^3^LD+P\[BM>c61ac8@A[0/b[-g>45BXQ0F;>UQ43P:5=MTD[U_SMFb[
E]4S2AK&/K4B+,A4<:B[;UJ\CSbU3VF,781_R:9MYYV?H1bT6O.UUEQ18;AQ=gQ5
OIJC+70QA4/R?P=5g5YO4f3\?\=Q[EQU>1I_U?HW.&3LO4I_=7BX3D2+GD(7=G^1
/O4BdS/D<bQH>NXC&Z9R>CCU]f1T=U#INVVg207]YVE.+)8EO_eO@fR\>gS/LY@;
OB0eV;28@(58/?HDBCM4#]-MVMdS&QILS#8#TU2K>V=cO<PU:R0DfX]9YJ>;E+Y#
(eRXA,_?@68,1)-bWRLC1-H_f5)Z<Y?K3.Je5#(_dYIWeUK^>gL=\)2_b<@+gT0,
b/Z1cFKO)+5c&36Fc->OaH-SHAB2LLV#UIZ<0g-gS-O/7>FeX^]RR-U0)CN>=S9f
1\I.8P2/^L@20c\9]W7VM20.UJ<CdD#;Z4,X,L-Hgc[H+C])X3H:(4;9g>\&:Pb@
8NX7^b&66c<&gXXML\,EL+Kd#S+JXK6K#(M^&R_Q8]Cd;N]5QDZRf.8DO&<e]WaC
^M,&OFV3[DPBdN[-,UdG0WWH:1fe-;-ab.W;ZGOWbNfI+9UB#BBRUbZ)))RO>7T3
5:d.[<g(OD48JX8Ja#0K159;[+WVD9I>QCWR,[#:3RdK&T9TgDJNO=eY:8VMTL^Q
9/QO=D;F(eP(5d5/?=7g=56K[8U.J/X+,BA2<5B.Q/I2[:4KSM1dYS&O#-2A36BM
/_(2>N-\&GWX;9PI<]VFg_e&2UX.F_8/_XQ11eYNY]BX^G@3W0BWb@4@cIW>]FR8
47>5\STD#D;d7R=SL(gTK<&E]fg&T)fFR<L;1aE7H_Y+CV=PXKFW,Fb9C<f1=V5e
]JO13\+Cc64WKa8aOA5;bN@ST>-Za&g:W7M&E=(V72,KMB<Ueaa/1LJ/9b(b<J,U
<^-C71,L/\+2;b_<FS+4F.CZ2[]^T54L6,dRGAU]F>G^e^Y__#W:1#4979?<J&/I
@)Wf>,[UF1L8ULO\0b)9486/3.XI=FEBFA0:<fdZ;^9N2U>aH9O/,]@0B:R#d3[Q
[=/dWT0MR]>3+4[daf]MeQ<DV@F^5([Af:[,0Q.KNFdREc0S1-E(29H^;Gc3A#<B
J+?>1J4d,HWMc2/a<-gLN>W;/W6<>.Ud49ZT<&B+2Xe^8N@dBBUD&TX5I?_KUSQL
#7<M>^S>),[1]AWYe/H6G=UUNQ54UZd8>GR^e.>Z8-^W=/_#Fc]dDMU(VKPfRE[A
X,[>E-3dYXf_02Og+ZXO9H(f,bQdM12_A5QDS1a#R(c#VbXF8?#)8[&>H?bbLQKL
6YL@SS#1\H.RNRDJOYKX)GS2gN8^_5T>U]8&ZIK/H]Yd_5SeHI:+]Y:RZ<A[aM\-
gV1fE+aNZ;Yfg9F=O#)N73XD1DaGNB=GWF)(&2dCH53PA&>:#F>TEYSaU&.9,/ga
DXB.OY.OX34Abe^3?(Ad5H=_9c>->V3DQXI&I(6X^ggA]_8T<L.c]5>?O/ba?/(b
U1b30JIV>b9IMSU-T]eRdWXS/Q=L7W),&d[+U\M4L_[YMLBD.5#Qa6;gO;.G/FUH
#1BFD\/R0XZCPPJ8093;@XDD2g>X3G_2LEJd6WQHE:J\QYFMW\Z<QbPV.^QTBR?5
Ke4[OS:LYf=V);EQWEgY,7?Ff,CUeFP7cS[E3gN-)D(>.<+HI^G-C<Q+G36<HJ]T
eU\4:IE+<.;MdNYaAegc[H;)]_6/)KIMF1>ScQ?_2f5B=(eV>B+7#<NL(^9RE:60
)XeBP7@9-H4@TNN0545eF4C@FX?VPZK3fI6L9)6M)F34/]a=QTC_(N/NVWR<TTCF
c98B&=@>4a6A]P(#)GdJb2O;\X33:Jg<Ja:d_G^_3T<N+M:G^JI19]HLN4MQ>4(/
6&B_#6MCD6]Ld+@1CDLE^BE95.(?K<_L+W[(2eSNdS^V1FaTfI.GOURQCfe\A/Xd
L\J98P[VRL>4OOM7\dO26H-NdK]_+K>d3.W\(Be5)a=82D[S>^2O^()4D4>MQ0^^
<3Na].7N>263:bXL/W_LR3gSL3:?#_E)?eG:Vg:5e2B-4HZ.4]IAM&/,M_9TM,dJ
e>OL2_9a_fJ9F7^&fA>WWN6be9E+>9d-]U>,Lg(>Z6bXe:D62XXW&e-JK>UbdZ)f
CM6T\8DOe^J@,6ZW+GB4Zd+JV+T2_gb#-?1H5[A7OU6U[,+C[K&)7L+fFMOLL0WE
F36U)CI>JV0Xd)_;+V8Y(84;Vb7ID-?Z(_4dN.-]79./V-MB/IKD]=W]Ug&<0\QZ
\<F<STKQMXZY2PKbQ+>M+39P_F6IB[&[[B+2b235;eK03Z8/TdNeEac#b);B9^2g
/?JB_C+U>2>Z3TD9L\Y0dSIBd@K_>9?A+NUS:VPD.8CC&IZR1LM4fVg9TfJ@,+d.
9HHQR+>_()W),/X@dGe\FcT:?X2UE.@dGDUK>IfEd0;B1A(6RH2)W3WVGOJ7@]_4
eBJ/A@ED#N>Q&^/b:\1d+0OHbK_Ca:M-Lb&10&Gc_U(M+f0?JHg5A<[?HNKYQ/c&
--L;^^9BXQOBMZ&SPSF</;SS))^Q5(()4dK&]&MQ0XY[&C?PG<[IZBZeRRH.M(b&
U]M_L-BVNF,D(V-?Y=P1dI.?DeA&SB1,a,+O?)O964SOR48dPVRV/,#U-BYL2d&[
)BWAYLDf<@J7GHfA\[.I-(O(^<]DT,PPG873W8#-5^,/#<3HB&,5MM;IEME5,e.Y
;W21BN>b&8fP50H7^HeUJg.P:\YW@RYc(ARgBX:XT)<46[9fI@:J\N+4]dR>^/IU
Ta?>2&-V8#H(BJ1-<=FX3/@>H-BY^@A--@JO8?AF8A(K[2JafOZ(^G17Xc<99_#a
U5WbN&M2YF#1/LKf&QI<d86,+><,UJD-O:T[/RDWefX\UP3R09JN,[&Y>0CNI7g<
F)VN(\R-1#9Ze@:]NHXDAFbc=X4N8[8K@H0>[X4/]<)-HF-[CCNN]cEW2=?I+c_b
H(8\&..HLBeL[1_.HPXNGASC_ZRONGdf9;=N_P&c9b,.9\#L/Y0IC\Z4[R0BK(-X
&(.ZaedK\S,+V1=JAD)[_fb<)P#;RF9@V4Re5DGEKe&]Q<KB:Q9c)O6M@LW(D\d&
Z)EFaQG_@XUN8BL2J8-SB)5&-2VSe-\Lf#Y=6-I>5:[L5)cb9K938dTQ2B8f\#3b
CJ]2a+7:N83S)_HMF.)\\Rd6;.,<AKU:c\RSFdB-Z9A9F^a>?2O#PGSc4FW18A]B
?&KL4?HHf2?1C#b\+GLI+#_#12MW<QU]<Q(g,>eKR;g>[[0CQEQ_Sd0F>[UF@OI)
EMH@X^a=Y_-GPW,U2B[FA>DZJ6D0K:^b.e#/(SH:>L=_?=a&K[R=6^H/JKC]N)),
GNSMVISL5V7PE1#@WSD\eB@0M;dJO5+P.B_&W5CWS-CN2,U=1TMOQ/Hcac;?e;(4
AY-Q06E.?<K2Yf);CVO^,PK^_dO7-NB:9d9N_dV8LYbeZUQ.63E0MdOg\@7c3+&O
^.?8_11W:+/6A3cbC50\V[6;E++TdHGR5bfIMVP.W1K-Z)eR)aERT<ET^.]Z]Wb3
(Icc>GBb=Y3N67H2/0(CJS&>MF]0:;-L5Ob\U(e+S:CO)9;OQ?:[AE+O5XD=BKF2
I-<]4XS@&EE24DP69Bd#(ObHgU(.F8<Y:EK3:9@OR_&<KWM;5C,eVd2V^V&b3L.@
R_8.CP\GI<,MVB>F(7QCF;&e1B0N+,N)&?DfYa6^V0Fa8/;RS(cYEHaZ,f0@)K_-
_16:[8+?K>3Q3\9@AP0<UU59C\b\/KNfW>GQ?gO1f]/#B9Q7RgT[a-3O&MbO#GL>
,#b6A1#<b/P_7.PY]b=L.SN)58AY@Y<d&f,7b>)((16G0@._6+aW9PgGB-7SbA9&
[7IeJTC>FGfb/H6cR9M^9R&Q)<KCbVPM\[\&[Mg-7M21FdT#[LR#Y&IT<B5C4c#P
PKUUc(L.<>HL3H&\L^D0>OI\)-?,RQR+JcOYOY6H-B1\&QTc6T8bGFG8VN-QO[V^
W1.91Y[;G6d4ANC3NaCTCAd@FNK+>dT/9Y-JE&GX>H,FXW<7(1BNYB-aD56ePc^,
EP4:N:,^LgA=3SZ>Dg=OM.bgPD/VNe.K-7+L<]&-4G]#F=01&;QK,#_35gBUe[S>
>ccS;,>/=W?gX5R([dEFMF[][X(0+1(C+L.V_:[K0\36JKL,_>6_6f:]5=6>0K5R
bgHYTW(G-=g6H6UAgHM533-@MbG:QbLC#<33?\PeQ]:6T_Ie1X:&+eb-:[cd6FPW
aBaC(G,RLVLO4M9AF9UG\IY]-AGHO0_ZH,>883.^X6aF(@KDJX1LUZ4/P7PFPd][
E_(]+c3:X/XL#QYJB06C_F>aSEc[/4_YO-/].J^XR0BH0Q^C@ZF1g]#3SVDG?+/6
e)#bcEKJ<F7XSK97H9E9a4:g5A1VY3GAZ4ZVMedVT3UUe=LS:?>4d007]-_:ea&^
O^?gcI)W>QFA^C]#9/+2O2B4(\5E6Ud@-J?221,]5A/I>WGD3&7Y<.C&DT:&eVN4
C1-(1HgDLY&[:dab+DfTMYJE,^eG2[GNaOKJ(.gfYU<.,J2<0fK?De\@Q9>)8PeF
RMY\0RAgg;AYZKd+89#5KH0]U[/J;&>(cM?R6b4:^&CT6dPD=eV1g[Ef]?MRF(E3
aN;5^KQ][g.e&U4UGTU)<P^caH(c0UO^,H0b@F)V7DOBE4^_QP5@(XF[+(Q^IJ]L
-eZ?&@FFAS1X7c2@f\Se^V7e1;^#K;cNb_eW&bB^+3.bLSMNFea5eXQ5\#fa[YH9
..8=P[FRcHcEH+M;4,54Gc/6FMM[GP:=HCBV>5)ObF59Bf(VSO)fW?F.W2+EGP\/
/;N)NI]_NIcKI(H)gO&N6(GFQK.VBg(JQPN\2GK&\[:JD6X4^^E<f;M>e4B;=G7H
2,ITbf]bPO3cG6ZMJMeD^a#2fRFY+)>6;gRC)/VZe14NN0-c:#Me9Z9Ob:.3HfHg
WF2X/dN^9cACZgTf>c8H_<OI7+,]7L&L91S5/fVdZeg<)/4+7((>79e77FAfgD8?
^2:1>fa3KGJa)2f@WGQXbc<9Qe]>3BbY\(UPSQWeU7:[TaX\M.W0eRC\/)V+ePX9
HI=8KS#^\=c3VZM1SP[B(a(M3NR92E-7GSZKcZ,AGKM^NJ;dA2TSP]:<7VNMF8_S
SO>a6>663a]@9FcJ,)NgM2:M[OY_2CZ)0[H0:-2HQ04YHAY5OEYacXLE?X[47L&g
&62UU3?;Y.T1=2_73@dG7LPgQa/17)2C@U1101HH-Z>;UE)S450D)D=S;>#Qc79=
(.QBTPM<?<^VVc:#@D/N91K&5S8F1I;N-e(Tc].;3W&;YSS#98)+,<3+:Y5D??WE
e;^8^1Oc)MQH4-+=:0>CSN+2gO[I5/4(a6@F[,HfT]A#?F-QWdN;K;C^.gGRRA6;
P+cQ_DbCWV,OENC::+5,5(a0\7G@1G+<AO[_JY;YQ=9DHSDY-&bE(g7@2MC9_O=(
PbSHJMMc<,g4I4]E4<PfTF/c:0.PJ/5-#9dZ/P73S-RH8K294K>+=g(OVZc[aU[,
X2P?)]=FEa8M++/LZV39e+(3V>bSZgUc\RG84]:deMZOg^^FP2;,aZH&FEX3g9;g
SS^dVWP&E<JQ_6d(g5eN6H60>>XN,.F3LcB7VGa:+N2Z&,.4:+2NZ)&A=V\,&QP>
WB:;M7K-U7e7\MaM&II8Nf:H6].\/[bc58U;Jg=1TUf]B3-+4>[QJ;@SENf13ePa
#DG)=9TFKNCZ_aZe(aO>@,)>C]+O5+YfYaO08=@@UE4L]_W&0M]F@YPb=DSK6Z=K
P9#cGHMCF@5,-daH<3CNWaW==(cM<BHS:AcWT/-V2(C(T)/?dSXGW?_Jg+bTH#-R
2A8b9H\.NASAAC#+RfF.&c=@;W_;=613F^BZS^:SI(O9:2E#^HUVU)FWfE.LdLXF
A,BYWc\=J:K2=N1J/.[@HI3T@f;5T0Y<]OOOTc2N-N,^_^ZG/?<VDWYP\b@\^)K1
db)^W0ec8B+SQGa2;6U8OO3+ZC]A8H:f0@C6,[W<<H()^Sc/?3K.VG2K;BO\A3?N
UOXYSf>88/#4,W<RfI&=<Z]&,8E8a)&4?[J5CLdII^_NB6IM1-E&\W],/LfRL2/6
BK[-<1W/(Z]5Z+B[XEN9ZcZ]-YQ[OSg_&,H:/1LFL=?:&E<^XZJZR]TW0<B7VB#<
-PcU;=4?5HVZNL+a3a?^L3)E1dO;W7]H\3dU6BFU/89eeS(LbHGDM.Q&LTIF(dEO
aFCNC)W-G/[_PD/\)QZ146^NVS?BMEW++<CFfd5[UBcKS105g)4MQ)XI#,BKLN4a
#O-3>Q;DK9faN@?33>A_)_=4=M=/^9K@O\bVg+]L<BSEAN7)SZ(Q;6KAY&_aH3]Q
MX=(ZGPZ7c[NXc@1b_EK>>IDZPTa1O[-X-TWbWO7_+11SJ#._e,DM0_;5#Q[;0)6
+4&,EIM,L9<U58_;eU477_:;,1U8TgB6Q&d;6bdd\UP>U@Df3.;Hc.C&VO^\ANaQ
=HTQ<+/Ue#FF?;P1S7\X@PJQ#EK=g]01N-3OIKKNH4PX1QXe+CSY&>1D(D2)D^@Y
4)4I\aAE:8+A9<6@;XaW9cd-W)9\g.S[G]/[d0H@MPa8d;#[/7P;L38VbYE<YcA3
X[RO,PT;IOe^Y67IRL(-=Yb^LPFc.UDeQ9K(-A21L,S&8ddYHK^C8;aDH2ZF/YY6
8&:ZE[gQUBIO.T28-__5T+bM0Z2(T7a2eR,Bb+\B82HA+=DA;4@/&;1(>;_TO&>1
^IL^XSG6UD;,fXC;(f3Q8S/F[2R;5.a8?L4;O,L_EbbbFPM/_/R,@FEBa&T#;V01
ABH#SOTRXU&e]])+[>N-S1B:H6D9/Ae&dV?AFbV-BM,2Q;Q[_O_(A,dZZ[@[B=JP
e,d]?RN@K/+cfGR+U)^Xa#U1=Se:30eJ,@Jg_ZTBfG]NDF(^U<KP80^A:4;;d7M-
)b867?[:/NQG^JaJ/eT?bYW=d?48d>#.a\FM]Cg:N46C]0)9M@b(f7GL\+PCUAQe
Pb,Ea1@_]BP[)B<fK[GU-)P61c?\V9bE;Sdf+XbQaOY[5eJ#J./FaH#Cd3OEIOZ>
\5QX\1<1KU_G>+LQK,\D>RIaDU(BUAR\bN+5cNUYT<36J34[G)PG42&):Q)3Jbb8
bY879[M?_7XA4Z]e8LBCEC5.]gSf#RRFPDA]I;cXWM#bCcf<7Tab^7BS#<gEHCf5
9Mf^><1f&(J?0g5&+D@D[MG;Fc4[>-F)T-=DK+VW-S2@I/fB5,+Le^BbCO^dg1]C
/#OA>3WQPGc@KS27O7&g0@09->)NRS&a5IEfOfH;f6IX1^fLWeE;=#)[Zc/CSRB<
C91XggB7IEIA11Fa#/[U:c<;DdBPR47-43J]K>58ZVCa/(0MaVPU)_BYU8YDV)BU
ZI?d/T9F>^>6(>W#\-bU#STf<A@[AHfVA?d.fS4,)YCW#6ZXUTda8e^:B0)b/5P&
8SSX]d,7:2._0?]M>2ZA6S-0W2:PBYa@FV6:MLT&>TCCe9cTTRb=(gW:dc]Q2_09
L=E:3cc6KG^A-UYZXcJ@O?d7Me/><&e[\<e+5D7[e<G@HWVCWZG7UV[cf-]HLVAO
gf57[;I0@Mb/X6^1^g,,URN?T0<aaA54]S3#<?C)a:3(,[L9/3??^-POg=T/f2UH
N8QW?eI@ZJcBA+Wc\&JQgP5V5EQ;:b)KdQb=Z5F?KXY>F(2^=+K.>MC^5&&OI\[C
^/J89UZ?C1gK=N0fg:Z2XSgBU9>T1/>O.<.L0\?D@\MWPZ;Z:eV()_-;A;Q?/-A>
XM81^771e(1VWd/3]G,6W8J-9dd8]YE@DCPBSTD/CJ?TDdb,X]D03Z1:R?Y0?4+f
_PM9HJ/POA37eB;L05,7G=dK,5f3VP.KNYADNF]>8-XE&&g;Y@ULB#C\(1>H)La1
cR=?.3;+.V^cGNXA\;U>>FP0;C[_b9)3?/J4:FI0].1AQ3XA-_PVD\]>=H]R[7F+
(]>&ZOIdTB0MW2UgCQ/8<UBN;Od4g)&0GfQf.WaAT;egB4YU,X[AaN.I8A.IUFbM
f1;f4=FCg=GBQ5ZDg779,O.,,.EbZK(_K9B#A6)20X+E)6Y4(5I::eV@@>4M?[7^
T7J=E5AJR+La([@0UAY_IJHcEbgG_ZUA=9H=DH3&^ee&_C.1I-XXGRA2YJ<.>J4D
cD9)D-2(\]Sa+\TT,;HL1/VF5\C4A8KHeHSRMgQTIAS[#SNPR&6KT<C,@1.IA9TS
QTNKV7?OYI(:=.,JHR#R<EVU.9)#Z,\7eTTcb0^Y&,[<eeU=CG-Y[0F.gTR4Ag(/
1.065SY^1;#8S.3KV,P:8O[0SAT4feN>\+WCZd57HbKfG2]]GbV=fMbKOOe8+9Q#
1;U&G@D62:g:FEOV[b8@ag&<aWC9P5>7Ie6\Ic\>4HN,H@^@gG5e37HfRFJ[e#4T
)2N.4cU(1O#9\b8.c.6gVVJ\g/VILgR7A3&()/-GB1AfQYXdWU?a33N4)M>5N0ZB
-NX-dQ+L2I\:f/5dZ5;J]Y>.7C]DX<fHKV/Xca\fBbKR_d#(?CY48fZQ)Z,0+-0N
^@)HNP2,P7,-:-77-Gg5\<;c]J^&MB^B[ER8=NLE-5W?:LVXXU&E0YAI/]gEC0;2
;J-g,<Td<KcA4BJ[5L&(^PVR)?5F:_NZRcaRQZP(#5d--a?PAB,U#&=ePS.TC^<g
AT_d,,6#4.8UNHc7DQT0Q,P,M>>bYMP6?G<V8X(3@]=&^52bL+3@#P@,^WS@2H+=
dgK7D;+>&-L^dRM6A<:>@H6b#DbQ3<70I_534JARO)>_-UU5d_0\Z]=5N&Y#@B=X
f.V0)XH2eGUBO)^dZ>d>(K;M:BFPS&[=IN:WaPCdTFIRHX<WbbKD)JXTe_fA6X?,
@\;[?_TZG.DSX4a)^B^9?,IZ;7=YM^>1T7KG8BG]N7#E)FD4=b4J_Y([HV7^b1I#
MKLQ8<eQ@aZ+\FDfOTULX\<gS.1b=FP6-G>.;J5?/;_JJZ#e1H\egKa0Y(;(I:46
fHa\.5LS7]#OJ>c(EQ[9;U],cF\d0.R,[PY(GCJ,[G?D9IIO2W&#2KHF;71GM9G3
bMW41?&BT;X>,9EFJKI.0-E,V,;WIPa;fSgGfJ=JGLVAM,5H(/[gO-^[IN#c8R=:
:dd3I0[-V-#A9_3&>_K[J<A)LJ2U[[dTYK<abNDd2Z^=3&F3G)Ef1+EV?c?N&Y\K
=,1B9:a6/^C[IS^,-;]d+6R_L>BYE75O(<2:cR0+FFF81V\2;E\FBA5[d8#9H7fb
fa1C2E6bdXN&DOX^/LD?gBJ(QC>S0.)63ASXA)CVC;?LEb=_-K1JDW.(G[-+4EJ_
e)09HVJ)^?O6aFO:SON0@_IS07+aH:MNAUSU(IZ,>8O0fGaCZX1O_/J);;eGJH@Q
,PC^T@\Y<0a7@)@>+P3MCK\(AZA0)5A_T&K[>[UIO(K/bVA:R<:;PT<Z&XMe4]b0
Oa-:,S.LYKO&6P/aP2_dD0J1>Q7>+?Xe77f\=TO,C<aI&Z(8^]b<PN/Jc+&R4350
;Q#WMgDI-#YF\WG0?>GgH<GE#LUF2S7I5&:=7@/?)6:HJL3QFDe\]6[.Ce/6A/OR
+87(f3+BY442>KILWgdZef#2g/7WD.Xg^OL^&ZHMZXYII)GHdW[KHCD7UdCHMXU6
/HQ#\abLdRaSRMa#67&dR[[;]WT9Z-NKA(JITYNgB[AW4H,&VT.M07>O(ceH<;)0
>,L;W>1Y4D?=)(1QU+=4S(\D;38c[WC7Jbe3(J;-__YV95[?J[V+Je=K0R98Q[_Y
M+D<bJf8A[Df7X<GIDVZBW;(^9e8f=2dPJEF@8<UF2Y,bZ&Y629Ld1U,2c.C63bG
[^3dG@)=>,2^&9_fD<24++CE13dQd=#EC1(5Nd5Q-M2T(,HB9VO+7J1;g[07X-2Q
dOMB4IE++QI?G(DT@5>\5ScKD02>Ab28H;GPL#?E:RE=&^a-ag6/G[#b_N=1GIB9
JW6+ZGSVR\GV5_QV:U97#fMLE.GaVb.3ZH/d^<8>KP>JQIGBbYD<VXZM2&\3YZ&+
C#88X;M:\<eJ9I.K>5,?S1;ffg4IgRI\Q0:^6F0da+OgB#fVZ2c8-T##8=Sg8K1,
-(BTSN#]LeYNT-YB7YGNfTV81-aRd.2bLEaW7G4/HBN3e<@9Fc.OSCO2716Z7WWB
Q)3KNG+K;USR=8OA6T9#(O+6PR+T?:A?;R>C\YNN3DC6a,Ub#7@?7JA@e6K2GWDD
_P3b<Z&Z_<#d=\)[6E1^K4S&]TQ04e[>?Q[bf8K,)0b9a:LU=S./[O,b&FY?2@P(
>YW[?R=#c]_SN\7XcEO@M]PDY.<KT;X;E#8VC+1U5,e_8VdH+WCITZ6T0<5/4\d@
36#4&I-I6f=<HTDC=.IH>G+d:AOLd:g)RE/:MM2.7O-bD2gF7^=OZON<Q<[_@L.f
@e.G&3d1BK9g3A&C:G6.H-LVWRH4cQe=YTIaWYUT9/[705V;EPI]5&:@,0_OKY[E
S(/VX.?B;4O)@+-F8;V[Qe2&^EZcKI,/@L(@+Y84DN+-&JP4RYF-6N=I:\+@-[(9
NBWY97.UOK>W(@<<E<3&IS7g6=V#?WLVa75+_e0R.0&25<JDJ2a46@&bXEAAIZQJ
&O+-7fA8a,36AfMH;]\gfS1]aaCYSXS,0UHbNVYQ]D?8aQcK\YQ)Z0GPe#LP7bQX
AYC4?DX8NHT/ab9JLXB_:1&Lb:)B3W0b,.+/@A(,K1dOG)Ze?5@@BJA/f<M;::N,
,WfHU9U2@=T,H-;,U]2N<,P]F2UHQ3B)-31)/=(N_0JQP-.8]NW^WYYEdR[HK>W=
G&6?WGGHG1.PJ4H;6>6KD\V<Ke.7AWJ\L85[]#:[+RBAP]8=CWC-ZQ,G^AEE/4??
./_f/^UM;Uf@B7&/5,UU[LDeS?(4<Z&;F&CFVDN9[_6-g/7M=RbK_?4;5\61?A4e
_N_Oa3\9NBa<(UMT=9U?SX1B@=RIW,-W4VW.:b^bH)F>V(8C.<BE=ZS\I4GDI:J4
FM@K(g2#7M>]3AKHJ/FUCARa>-B8)5KA@e^G)eH-eFHPge\\aXX]b;5UR[G.B0DJ
ONCJ7N<EIP>#QQTEK+H073^aEfG9EWcUec9G,Ad/(9T7ZMfC4aK#_F=:ID13O8S3
G1ZD[GH6E60--(E<6QRVJ?L]LSHGWeAC8[H@P6_=GZ;F1;cA2^PMKI<KPME]?4<-
6b9UC+c]J/=:M<g6=#@C53HW.]B:dJ;TVKGT]HPB?#(D[E6[IJR3=TZb=U-S/83U
M(9D<<FWf)MK1R-T;bPXORc&f(##))DF]_85S944UKXZ_:Z-,,<9#TQ@B[F:Ue:F
;E&ZX5M/.IY..cC\0T=H0B&P<RY[J(Ng/7\=IPKCCP5Q>OWO,_)7H,aV(+@Ie9gd
82c2&&&CaG77GBY^.V,NVbGJ^25E_4=14T)VED4a\?Z]#5SBLY-@9I,H=CT0)Pc=
Cg0E:B9=.-EE.\)8+#)V)F3)gJUXdO#F+J8LN^;U3\cUUA0CI8?HQ;3>\TdX].<T
TPg_b_#XeYBcI^dRZ88,?U/\VA?EAQLPD^=F/VA4^,2Qcad#_R8>SSU6e,X1+e8^
X]LAH.?eQX(:B9[;Be/;_(^MaKAG(53P.N8#Ie^]>_1)7);c#,0O-Lg6g^8((,dM
>E?SF(#2,[dYgX<:JS/L?:JG-R:R-MP3J\VeIM/>X?PD/?d4,\=YS1d9KQYD\\7g
O[e?US&g:eVO#X-CVL0^Z><]BGX.W4./:ZfUFDTPd-CG@_.dSaG295g_,>HZ/L[Y
)eBNAe-RY>N/9[];XFcAcbg3@C>&9/VbC.d5XQ\YC3-X5]UK1Y/e50@0DE7GS.FB
,W@?cK,)GL&I3:GNCe+b>^Ua3\PM6D,=.NR9[;^@YNDNJ<UX?[Ue_#e/Y?BD,eXY
RDL6bfB><]T,&Za(dJ<P<&[6<f\31Wa,J8T\JC6ZD7[((@WNIB:K@#U@4cML8K]A
N2A0P.:AT6X^B+YVMRAJe^F2VZ<c/GC6NX?UaLZ&-;bWQ,_1RbNeN=M[T#,YbXN[
@-@YD^]\GA=P<OKHBb(T+)352LG1QHN0Yff/0D.EK:a56b3P5<:74DcX(EgEBcQR
W+#/]3UcgTf2ZC=@S9cC.f71a&Q4,Rf7dPWN7TNZJ@G?AJaK11<SYa/dMPYbdNMA
aGJ,08a8/FRd9cQ9,LUO4BWY1:H16DaUI]4<MZ0SG0VQ(P568T?[9E-)9GZK=FOd
=YB:J8I++V&_cSYMDYUM-c:(YTbC:,bE7DH-,D1dT/V8+<B27L^\.FA10PR(2OfP
>/X<GL9L1FeK#;YOb&Hc3D)CPKeQbeI?G)-^-\8JILJ[^_@56OY(V-@[#:RU5L/e
eg>854M>fY,Q3&,FeT=FBE5b@,?=I<Y;Kb]NW8?U>Ma=IV#XcF75c[NOU41PPN:B
dS?e=YQGac0;E1;F-cB5.&&15XIQNAS_\LNbNfEASRF9XZZLPK6D@(J]f+)G_e7g
4.):K=/:<eNfVf\6&FW1V=R)U_6dZ<HA73VgE>KFbY8SM\gG^Ee6IBT:A]]cABX1
]TD8Q^eW(dY^-KSTO@HV3A1M:HfJ;\KJQW)OR3[;]+;c3)TbVS=RA71AFVAP)&FU
2RVf>6?O#Y;2CHTAfBFLa?bd]#A&Fb#Z2IX#F<\9/Z4MDXR&[P7#045.bB+L9YYI
9/K2N7@#+_9XLc4+COG,XgZC0=4M4RfQ/&?,^E;]]S>GBJ+S)4f6^D.A:5b\<7H)
_0M?3MOAJ7@fZ.a@Zc&#U,XN6RI=2Tb+WD+7[P_e)SA.S/DJ3K2S53He\&VVA>/+
A/I@b2FR6e3^/E[HOe@H#3eK+H+f_,d/#5T)/XYbO4K<DC[N\bd73&g1Q)PQCY:#
JD@9C;bT3I[O&gH69f\()BK5>XecV99PS_,cU?6Y?UPWU./e]TQ&MgJcXYdIQe4g
XJ<W;BVY2[,_IN;_XH.;NGT?\&OS7;]gV4>V\->&LAGX>2/1JdY=UAU:<H>-&VI?
:TZ.OORKSE(^3TOd?@K7GIaT6I6f<2,=b,gPa:475V7OeHHF89eKG#8399acJ:#M
\QATAT-V5HVG-;1,SC<6[Bb5#9B6c9dS8=S+BY_91@NeVFE/J78]M7.V7LMD4NGA
FZe??\9UF;ERJNJAX;g8c/Kd(WbB/O(&I=_N37EC:U_eaGI^e5?.ZNOA3;3@:8DJ
,VRffJL0=?>COG#@-7)V6gK;+cQ9P(RL7^22Q@CMGNH?<_bDTa9@g)3^E8?Ug9>Q
4Hb1WIT6b0>_eSJS]PZJ]c&\R_IGJ^g,HMf9;QVD2:P/W#A=NMJ]cHRdS((T>B[B
<W2=B>?1eb/6D15OeJ^?b4X_dQbC.P0SI9)UYAOZS[TG^=bO:[f^cgTSD0TXA7Xc
4-Xd[L,=>PZ3/gA5MJC<gS(D1.cb?Yd&UFRRg2WRO3F#\#:2;C2@^MNX,3=B:5HZ
4CLF9K\gY\0T71<ENPe.\3^KUN3,:g)eLD4-(gg9?#aIH30=M<H;28REf1?:BH4J
U&5f[V(#(?ERD],F3AY[f.UQK)M4;9&McZff0<>ZJ1^GRY;3C(@e2AZ36^^/8S,4
Hf_fOFJ-.7UD<GYPeY6[U,BFJR66F]^GGg7I=/QV>6Rc4U<fGfCOIZ_5M8[(H3=b
7+5(c4g_:_<@ccW.:A77@Z?MdJ])_LfFfJ?P2.#IN3c^I\W0GCXW^f1,f-.[>-QC
W\U.cGT5^&GIc4=KG0Na^PgBRN);(+30;(JDW^Y&=AC&I5H]aU\_T+Kc5(@7XWa=
=[,?U&5>Bd\CL[OdQ2dV:f8&WBa@N(_6Za(>J^b5fPSgH((639.<++>Q:WL)@aVc
SYLOJ@O1DE81&O3bCUH:g(2,ULF7?,.GE]RZDOAJ>31^6655G?C-;-g\E@)RC1<b
KbY#dQC(DXM/.Q/:BTaY.MMa3/0B^JG051^QLZ:[g;KDfX6IGQ9W.3c3)AaP?M78
aI(fV,/e.J?/[HcX.cW=4Dc4F1N1g^?,:-<Jc81DLKDIa4+HR@;=?KQd5;RBVC=c
5gN;YSC<fBGNZL?6+>.P]XWE0?DbUUe(6W4I<1cC;_U5cW@4Z#:KH+J<(S6H#+aQ
MTB2d<2eRHg?VJ/+\+\bJ)A?L^-[UZ<b3/A9GYB+V^L4[KJ+RG;Ha>MIT(BgY@/d
U,@9/Pd3I92Y=?ZgSM4ETSIAQ-U,@B(,B>cgcCd0D;,72B#>Ka=Z-/b@Za-[1A)D
]ZbM\+:,KX<TM=(2?W(c6XabEe;.XMY(#d;O^YAOg9,5[b@#AXYf(4H^<a4Xd(Bd
=DAAC^fYE4S@]KObE/U;C?5^T=WgQ?DOd1c@a63Q6BT[J.(BcPP4QS-J5:V#&ZS[
JA(=X4.F3e;9bZI>ZC)NVQDc[]N^&_eNBK)/2_Q\AQ-b^Cg3=2FX/73Y8dNZf<?W
H5N^d/VRPR-[5#VKJ??W.9:Md=O3W]-?G=>g::Y^3fbV&BeN)U39A?7,.YR)\I2[
55&@/IJX]3aL]5V@Yf:cNF1WTXV8)M5+U8KWFNJ1@>NWH#F7(X@fIABb3.E.Z1T<
Mf^W[cRA=4@QC^R[AbVL)<LJ8BDY8SR/8B3/\3Q(?7?63R(Z>LGeFQ:ggbLZHc7-
#-U6H93?)Me\f(?^EOC61FRf#=LSEB_HYHS)WK]L)C+]a>&NED1bfRFLLK#cYMN6
,^NC4ce)Y2V9)aD9C.Ua2=))T)6KNOAJ1AF;.T<)_][dFAR#EQ5=QW-K5T,&UO00
@B3(I[H6F@,T2LHNB+AS-^T3,U@a)Pb/X0MGe5MFKd6&1Z_NK6ZV9\,DJ5Y:QW2-
O/:=HA;ZH4a^RdZ#@1W[AA=B6CQ.1RUVeaI@I^=#b??Wc>:8f;FB>-K)b5H.46>g
WSXA^)[#<gd:9(KdS/CEH_U-5E\J^/1gf)?dg(d&S,8)&4Tf6b]1GJBad8g:0Yb>
N2gBgccV)LSCK,&#C:]DS9W2ab7AC9>fKI\c53O3RGZFYLUGBEeI&19D2:85aEf(
.fP?^6:B5E.T-^<gcc.TO\9c1(E\I)Z6H\?4e]2+<[@P2=+d40(_cNXY]SK=M3ed
/e3H4;3]bfe^K2?(EO74abOBN7M:-bX;1?\7U0BZX^YXI8g=GK/N-ZSN?F.+UITe
F?7ZD<GF.YYY=Y67Ac>7&(cbTGVD<IS)+;5)(4?8/R[33E_M&:4KcdJMS0M<C+-[
5RGR:b<5F2)=Y)c3+?J))?L88b\TT:.bg_ZK3V@M#7A9XTVK4=9P=f78:82#TJY:
AA6PZQ#WU+W==&HUe#:=7ZUSS+ffPDWG9[6(aPC,@cG.,+E,9442D2M_S&;5VOYd
C(L3Hc9##8U&6AO(Z::6J=0^bH<c1Q:1d^;2UN59eCPC[51KYD[P0JIaGf>W>UER
_=>#cCX62GRR(f(+g[4T-)C.cdQI])28,8DX_fRH96GfPA#-2^Kd(Qgb)-NRd^C0
M@8I;S,/W_.e,/QV<a[IED[.X3U/0;5^>gO:TODR>,gfL)4AT?846c#[ZTgbb3P#
_:?5GTSP--4EDO6^:5b^:Ze.gBMC@&]]&GX[_V0=+T+JcT?/C+A^+-a-U2:=cQ[M
a2e)VeH\:__F.G/0,-;Z29+fMZEW9DIRCHW/(c:b(+g^T.e]eX:.L[W&\b=HFZ:C
\>G[PCS67[;U(Aa;?V2T;c.6VH24;E)BG,9=]O@NU6cMX+#5J0(.N(&&\UGbg(gX
f4PGZ:#UM;61@]+KagH\FfJ<TF.54-\1N?Q/N(:L69fI(Qc(M_KKb\<2B>BeZ=F<
RJKS4-e2_1Td/,G/09fUI5&38VUK^=^Q:5OOXdFYc[fNR2\?Y8YKH98,TJFG&G81
PW+(7<PNV@^E>D?G.+(E_aP:I2]QV/8+&8f<>M<8.YS9+b.Z^HUM<P1T:K516_YH
)+aH>1e-NQaIdE[;ZZ[.<_7]2^WD/=B;ZPc&#9&DN8#b8/U+K_^Z-44Y@WX2c:SE
6dQ2=+.A4,#9OeEcP/-f]1XI)^J(Zf>(7\ET^H:NZ+2Gc8IHOP@>2BeK-AGM9;fO
9#]?aSe2P8c<gQ#f2O<?<KDR,&W9X,MEf4a:=d?[PGWV/4<a?I[9]87ZKdQDFH#L
gcPbQ1]1BAVZTYgR[b.)CBS=M5P651_[9ER1A?Z_=]+QJKA[VOG#V:89JV(R12aD
f:I3M[YN4#6-M;;-3VKKGTK3WV+GHHNeW)QPC+/E\2eX0056M=_U^U3>E3;Z7d;a
#DA\f\F4:Ag\IA,bJfP#]DH[bK_#6,^T06#WV7gLH>_.:#_<c_dBS[0+9;CI])\Z
>TdJA&-UD_#:U(3g#L&/DY8G4d[TcQY,RU:;5g?7EI0c6\;>#3&gc[_-]4YLXW-f
ZZ]HENc^H4^cc^.-f:K-MB(.@\MXd(Q\_OI:.&P8CUE>RbbPfBC]><\cLb(d2BA@
=R]d((ETLRNLRL]UYJ@RMY09JJXKRV&O1)HDVM-c1;D80Z=R/J0/V;f_X[&,C.GZ
>(3dHE^;8g^7,\#gCQ<,X5A\#)2@Ub=@9[ZZ=+Dce[14<-A[F+Y:3.11ZERFEXST
0/-:_UQT>J\GT\43F/f,BS=X_b17<eV58QCPS_K2>/FeGfLB:WJ?-TD==Z&4<=4N
9Q?3b;Y9<R75aF4+R<;0AD0-E.4RO3(YfWWI5OBFeEQ[^?LI7E2#bB13EU^bZf;7
f:0G-)f>SEBUD\DfOEA\Gac@@H/V#HIAZ[cEC-H70=88AY?QT8IfQ]gX.>FRdMV(
Z<aMWF0E@77RL8PSC6VaH<>+gV&2PT_]SJ-b<LJ_(+R[8(<aY2]R)=[c2T7I=L^[
=)=O_9+V66CK()dJ-AHR4=Q#O9.IMMQ_cMd_T++1GdbYD,7;c@/RL1=-:J\//VI:
URB-^8(cgUg[CLYd]IVI8<KW[RfB[?8-O&.)5]-9gM3AMMF9<N86=T4]^MG1[IAf
Y+Ke/LT&<T4bZceA[4Z=@/&VAH6)fU6:VTTVRK-VY=UBA5]ZA1#>:N+X_eA9-/V9
R>:[Gd_92AS+VR]X8N0U3ZQ2VJ&g,_T(E+Q&Cf3<0^]?\g81\:@K@BR]IZ_@;JD+
SLf&P]Xa_D09&O^4.C:2&=8B[>32MY5fdV+b((N@C0KS=F4_GdZTgQ.(^..V)RXa
@c<4MMK/1_/f)Rf<[=XbSE_R9?RHE[JUCU5A:8^5OUa_-_g@@Q3BF+=V#90/UdYK
\VSQ2U/=g_^/fIK8SV/#&,VB(b43RJ1XRCQ24T8I#4:;@&&C;[X#MGfU?<8@BR&E
fZB>B@E(I8PAD@&:X(@VbCKOe\5J2AVLJ&Wa-GLDQ=KT4P0YS<EIFV8^D3faT(J>
V3:.1acI34BRA64gBGb:6?,V:LB8\dT>OR7)LCf\FTZ^OXD@OT\H^)16+?#10BYR
Q[1B\IFC4K_2HYb.4AQ;)B9HIP&V>HD7a0_1OfbRBE&,?.2G[#f^>:KAbFMWS.C_
_)&?&Z[8H=4-BQ0;dU3&7BF+-D[3Ye2?&QV]d-_Ta+6>_DM@-)+PB_M74-C9N4gH
+_8[RAQW;_N>)a.TI&S=,9:]7U9SG8BQ+7OG\gIdFK+C=Z_=WD=5V-4(#\Q-&)EX
6O7.V>AX853#V)LX#eDLOOSa4FVFH+FIDUJ78Qd5?VMGaT&I\>UND6d761Fb(19:
3JWS+;/D)L,g#^EL?L#1+BY(_#4F=fE[.R0.LH19E6C=1BggS/<e,TXW<+;DFB9M
G3U[A:8Aga4O>J=gL+IXa=N8ea@bLfO]N_RH3eMR/5\@B^^fP&(O;V<\=(?\GRa_
eVd]WFHWXe#U]&:=dM7W]L?UBNQJ#d:6CGZ9--P7eO_1fXJ_:\[e[08eEA]\X9W1
.BN-0\#cL257@86/7I@5;5PUPW/\c5fJ8YC-\1gYS7?ALS3M4-<IV>E2:P#_R8.K
)FF>\(Z7@e-NO>>J[7G2YF]5(5T&35.4bX[+\)6G@YbOe?ag75_CZJbWKXK_&ePV
9gIBA59R424c00__4bbK1B^UD(1:[eIQ?dHXIT+>:(Y/#EWNRZAN\O7[R>4WVe2J
](F8O<L0##M96NTAK^93DUH_eBD]8143\ON(8gUFF>@^L]A]/+\_9.X(W@f(a+(Z
P1>Ug&#W>D>B-V4Dc)HOM<?B\JbB(H0TD1L5O>5&_+YQOQgA44g&[f_dK;AfGG.-
>ZLZP;9#TI(QCU?f=c25)YEKOdaO>C_^=V?\f-&cgdUB\Md/e_]8aggWQTPJ7_8f
X#[G]+aB^B/EA_G@HQD)D/OK9Zc]]1fWLMV\]D]L3Of6TM<;,=V[;><Sc2ACM(RK
D/SdeS9.K64.)bf+^&L,V9UZP(E(T\0Jb58HbY3G(E/Y2/gFCKAGfZ(5X9K&LaN0
TgI?,USKfdVL(C^6?5I@[D>1UeJ@KQd&DG9Dc/]1>D4:>(:_(f:gO02TYGWa6H60
LCNa+b_UKN8K^-3COR7O,/14,(f7L/60N6If=^g8.P6[)DENF48[ZgSDO/8LaZU.
I-f<8;cN9L2YgT;@f<dMRPL6=?,0:SW+\NFa]GMFCFLVXT],:A&R#1@VKIZ5+g?0
,=:7XdB?dFAS@ERG,Z:-d[fU[BEe>[VI83RSAfOE]RY@M4>&#&-@S[Xc-EAgJ=K+
(Z_.)HZPF3^,FVBS81.QI#D[Iag<#//&KTJNGIO5@LI=^K/2&8K?32)Wb6+W+X^0
cV9^B\E8U\KUIGZ0[VfB[>^&S._.ST9F@gG>.US98:SL52IDJ<^M^X-bI>-@W:e4
a+SAK\df(8LR(R/d>4G3Gc+efEZY\Z&gO@OXcb&HR:\_#c9@[UVE7d8A8KRUYfe]
2B<8Lc.4-fZR(B>.C.9D_d6NdeJ-WeJ:P77N+6L#Y:aSA1&4?BVN[EbKI3Z@F)eA
)_IeJQ.S3LFe4?]<5ZE\B>1BXEN2,\H\=503C8ES/d#=>V48^):XZ@,72>BCaf9N
C2&+L3??D+3D:IAM_?FAeK@A=:O]P#E/a^7VA=TVdKV,+((.I0dH(7d&cS&f=Z->
G6HTD?V&W)VN,L@LV2TPcACcI1.e<8baVOC:dJ2\V3N^TGVIS<7Y[ag86/CX0FLL
E+U)Y0H[S2T(P0+:;ILRDY2GSHJTRI:?5G,f_+O=&e\)H.]BJ:SIOcI8JB2SYEK8
.RP?ZPK5;#=]d7eJ\/5?M#X?&089[-R0H)NJe;K&D1dCI6B_DF39_G??]V?#P#>^
?T[G>R?e(6SE9:^Y/L72.,=)H0]]LOL_)1GD5-PZ?P;/)VMQ&U0_2G]DVQ/4G(OG
?BB&E?W9&7&5<\7B87feA(SN-<>caMV)ON,-PVL4>U<6aYC,WL,0GA1D\GcB72bc
((]#=>2Y2APPFaZW=aW\U?S@_&]L/R.9<,K)7S.;Sa?U/]gR?J\G\+g+(eZ-5B06
g@3X(-F.P:=S8I14813^KdPSKZ>+&+5<L0[P&_b8&V<0N#5F3,H3<02S]Y#==0^@
SZ7R79?V-.7=9BWXDO^10>.>PZc3FJ^UM4H>XCcAQ7JT;SOgS4ZVD1#2[-TO@5J?
6f/T)I<SIA0G+N<=(d2N;,IGI(c(GH8EE?.MEUJ8Ma1RI_0SHHfVU[X0T;P>:Ze>
)dKddZEV2X#4B2=0+KVOfH\B=e\5Z?#EBQETUAJ^.=(P.a3+EP2_N0?gNQ50HORO
.Ec]PKaJ4=2?#P@E3B_cU7#O(,0f)95PbE[/(#ZD3eGDNR78eR7QbT\JLKW@KRBC
MY+QC];[<FI(=->4R81B?,NFc,c5_AM/@#Jd#=6J#6YJfQ@@-SHF\(=HI:4J#dYa
GW:H[_HHMf9>dK.@?(/]fZ40:(fI6I9HG;#+<-KE)7BXM6a8e;ZP(\>-B+a@8E.<
6=&?\4411ZDSANaB8:[21[5X>T2U6=a=>=fO/5U)\7VbQ,4IR>f=<^6\,)H:S_L7
YFX\C6?8&dW7g#E39>@#M2[UY&-:,W6:IQ[cB5SU98__e.G)Xe6)OHY[1&618,3L
cI;XJ=,+007ba(DU&O,D2>\1HR03e?]H9(g=,(V/VD+.AcJSN2dBcV<Y9&Af,(H/
2WINRgIOF-9NK]2.0:P]07-1[QEa-,BfJNe;d[49c_>V=)N1P:cI@?SC[>5B?SWQ
P\DE@Y-?2DGT+1[P+I:GI(,;6F8S9BC9]MJ=/aTCLfWET64=.;EW0.c&Zb-,_^V#
RK#)cPN8#O5MR4>>Vb5?BfTV]H8J@0PA#3OVf@.U(A2CB-dI]OFH:-Z3/f<d094B
SfK3@_S43-<(5.Uba=17#9&3NSZA<:]33P8VUO:HQDKe#ZAf,O,@?F_ed,M0Q5^G
UAXF=];T,#XN90<,9J\;3OeJA?CP^R17feD?H_L9aD]WDea(;S=VAA(77]HG-K6a
5G+6+6E=C-8Xd=C>/>0XHCT6<8@<S((e;/[deR[OBG\BgFS-.Y6]IaLGNaR2J445
AO;3^Q\\5UTAaG3bFELTC:_8^G24dS?&N=c6NMM3\J]U6MHG?54[c:A[;_,U\dd>
=9H\SZ@U#&(Z8OB^^Q,.1QOH<+NFSPQI[<[[9\]OZ#^Mf@_O6(7Z?ZS402<YR56.
X6ZXMbKO3,,K0/(Q]A//QgI?U6B[Z47ESJaSU-8cdANBEF1a79;MFb4bS;J];[K1
15^Z:dB-]^22=PdG\TVE^E^D-TTJ5OL#8R0&&3C(MI+I4SM+2B6,-)RG9e,^1B\C
/PVZVd6Zc<fIJ2M@)-H&NCBOMK<YP1+1eU,eLSD&/d&NLF4BcbK[157A/E=eWX^;
cYLSVF?W7\XPAYI^9?J:bI#[Ue/]S.8OLgIc?JQM(B.@[5HfW6QJRBUZG8CCJG3U
bWEK@SY25b-24TY>2;#S\Fda0/=KRAS@(aA6+9?>8d7O(:SMX[b>\WX0ZTPYI^7G
:1f)@ea4S[N)=&RV16E,c&<QSW3f:VY0)U1X<QY,W,/)cdYP#OP-JM#d?a9=:Z^<
3+E-39Wf]TSR1EJ^@<?;A+@c-(]67/C<B:9\eHRacK>1_H(W4Xg7OL-A;AF#2L9-
eU\RO>fcA_a.4@fMeRb165S/GWP]ce>VL&WH]7.UYcPX9Xf3c-e.E8Z\K\2d<#8[
)/6BO?YF]K+EcY,2[?-4JA5+S.R]fP=[&M11ddgG]K7#DFU6F^&M?D,__(eZ/d1I
d^AXPY;876KICOY[15Dc-4ZA8DdUG?RcB\Yc1A<&)8>RO1L;g[X1;N6;b16MI\J[
-P9+,)L6:eAE=[19VfL4+S@L&+\0[cBDZT)JGRZNUc,0OWD@fR--K6R8,6^<GK\&
\e1WQ3Bg,A+?RFGP6:MVa(UeH[F;G(6LBD(\-g6<?5.ZL8OO[V/g^:Z4A)8]?<LQ
&/5B03&AW(Y.^BEW2Ub@R;@X<-T0Z)DId&,?I\@&-O.gV05Pd;[/S8>OC;NdT@<^
.OU:YSNO>e-aX9F39[DdJ=BD5[H]RX=DUMH5.g:SQ[.cF9NHa2fc4#0O?1Ta0QC4
35[:-L+WAe8S4G5NZPf/dT8IedRDd.(893E?27T@ZfA2_F9V.C<(:+eEPU:d9PUe
fdJ7Y,\W[gF_cOCY9f)7<9>ET-G-.-5&NJ?F1+M:+@\<6Wgb_Me^3<A.<9I_HXAR
Y+b]=Sd?DWRF^ZMFQ+c;.IG-^KP_;LdOIVHf,AA#H<@g8??Kd]48B[M:8[5XCFK4
Tc8BZ>IBeT;0:[UVcB1M0X<Cf6AD<Z/69P\#Y8a=N-039UY1.2UYVX1egY0J(-MY
EK?24NR-Kc+/D6\I]ICS(;B]KP)VXT50W1-fe9eNc[P2_?33?JH-:3GFbR>\U4>M
^[X_1(7-g9/R4J;c;(5Q7J3(KJ#[/+P^IQ5\J-K?RSeD,K,@QB-7,1LgXD&&-G87
[EH>bgCOeg.WOC&EZ\S7BTe@:1#&#1V4Le^dV(2#Ge8Y6(N>1cJBXa[5HNI=B&G/
efV#35dFQGRUC-::/?T6K/-HK,@]g#9D@eHe9cHg[0?IQ.X[HQR.&3gA)W)+<)RP
Ca?+CZU7L(g2ZHf\3TIPQQ&9PX_N(;-7PHPg8<dZ>U>JaVG/,8T/A)H^JWNaNg+5
MN==>MHK.,N36.[2<R+)E@d2/e=AUV:=eE[WO3O)JVRW=DZMS05M-P8U,#)6eD_P
[M\2DK=)aR_/W>/UJXO>T,P;^FP>0JQ?V);U@-UWBMB(PcEKeR&P\&XL9B#^c,6=
G?PD@a?Ra2_Pf^]fLBV=>ML\2IdgR(=ZS6c+#C0efg^X;5]-X[+POI/\W,)e]D;G
S6eZ32EV.e&R#[OQR(SL;V/66G(^gBPL2)Tg;S9,4;WCD9FN\ZZ2VZ<#5Q_/9S_R
)>J\4WZM?0;9dVKX(((TR)N]@H7Xf.D2_X-Y+U95?3eQa,T7K\7PL1&[J8#H9[=6
M;,A=e#:GHCcHd.@DIXSCFPA^7d4@W@/b-#CPTCZ6QTIKXK_fFX+B.&L[(.K]-U^
_UdK2,_H#PL.C^DQ^\+W?1(Ob,gLG\C8BfDBDaQKYgE/@)P&P0@4R>U19(cG^]@R
a6+U<PAJ]dKNI.AEN^QQP[/?D,egB06+LX5B7CKK.1QNCg(/\)-RgM,X?8EcR]&6
1+<eCQTEKY0C-Q+(<RWP6g2DRK_WJ-D=C0BJ=/S/Y&LRAU.,SVaPN1\5@?[N<]&E
6(4,DWE:T?KcL<R4<Q9g<&YR@3Y#g5681;JQA^A4b9V79Q_H)g3SOIA3+8&(CPDM
N-cgC;OF&<L9R05]3RIg^-cCOSdK@_&8aBSM9NN&De_^I)1JDPL6gb:J(F1Y\OOX
bNQLR=YKd<gAf&>?-e\D)gBUJM2Ze/>KW6L>3[=Q6G)O=U_f-<DfX+a#aBgA#NG[
?JG;.#F8:cP9]UH6,=84^,DddCLL.@;VIJKS#WY6[M=3/Y6<F<>Z57WPNGBC[IBK
LH80WP8&D+A]03OB)Hd13[Y=O3^<a>b^>0C:3@Y=XY:Xdd>,#0E<[=YR895F;HG6
gY(8&Ab^+77[R35d&IWOXD;A8OT,TSV#^/<.fScW]bSb\bB:<LQSgd@5]^E-XN>N
J=?358RT2=Rf1NJLRFAgWG>c)-:@><P\>CP^;FDGA)L<(]b7D=+DN/e>I&]S^V\2
7NRG,egX1^G&:WAdR4BSFHCY0D&(+EC>589e]=G@HO(A0LK&6(a_7WB@&e/S\>@N
ea4X[WJZA5+3#@1?KK#V[K+eH.GH5C8c5EO=U7^:8)_W/@#Ug1<L&29A#1\I)]dG
X.+47;@P^[Y-d@]HIC>M7>&;:Q#e_;AM-CcXe_5I849RNf#C]S^aH9+VURg@UVY[
AM;\P+1DDdX8PT(.)T+GfKgA?;<).&Ad:GT1\>bL4EA-g([4<:W]c3SE0<^3UAMW
fHX0]FL_BBBa6VLaCX2daK]Q=RcR<0f0:&gGD6JN23;4=>1PbD:KOHAR;^5WCeJ?
77BD9U)3SU78J[F^c\VYDcL#I&32L>a,&W_4#@bCKeJ86USM>0N<BV3gN;TFc.NO
BX+2eQRCZN?a,CIOV?B3.KWV:^V=Y&eXAINQ<KX03_?AO._=08e=eTPddQYM6L)Y
527aM1V?@Z-701ZA>eKQT<]aVd>06GLd+N(>:<1T6,9&V]H@831MYG/F36CZL6S5
&V<3FMF4UUVdUH-KF=5;I9[_M[X+[YQ>c;@J6Kf0fF8=f5gA.gc^Y(S403+;1L2a
cD;>;8\TgP=CS7Dg-^A^,FG89O>],[E_6OYReYdIW22I^]K4.;+4gV8;QC#0VY<b
1HbVLYF<dM?AR##?EdK(S,A+.[=cdU>3J=FCPTG9P.Wb<9C1DBK/fdfLcB:0[9:-
Q<.>8SV,PQS;,^c4DN(\VeZ@G^\#8;fEOg<RX[V^I6cFfS(\bf[6Wf(GNG@8^PJ?
H<K@a<V45X?OK\OT;JZ<98VP>g@:U&N-d?gDF)eZV:1UD5#H,Mf6JB9bB<ETZH<K
.KM=d4WM)/.6R\9##S_.BCfPLE^+0&:2R[W7(NWR;11@cF^a=^QK80_88.R6].&B
R>5X.T\J@/&.]+4?JEPNA#M4=:S2)5O?N5+8F]b+e8Rd7R#Y0=E53,4><N&AKW@S
Q/7,a7fcEL[#3JeFO[R>1O[[5&1O.M[@Ga:3EN2M[57[/aJVc8S;2[3,Q1.]QXf[
??@X.WPTQKabY_FMP:0YeG9Z-,109DM6/:;.-WXY1H>?(AeH,&A)0^U#>cZ-Of[?
>-9BbZ\(fTH6HcJ8:(ZESfc\RJ8/0R;F0ZfH\G,20Y:97\@9_K\Cb^:\@g2BAN,C
S6M7bU)GIH:)Y4g\7IUI:^;T>T),XGQ+fTLD5ZYPQJ@L=f^ZZF<Nf&b=2;MZ:YeK
AZcaH6VdU-SJ36dEK.Q31.5.c.Ya^,J1_[WVA#U@]M(gF^FdW[;2\O73AL<S?V4H
)4J5B/[?@-P>=WZ-FZ&ZF33Y\,SBe4=;5DHY+&BOLMbC\F(bI]IPa)PZ571J<?P>
9:0&34XVgK45_[)(3c7G\UMOZYPR^aQ9F380;21?2c]FWR,6G9876P@R0T<@T[\/
B,X406P=d3eC,N=BcdCFX=KCeKYEATD61dc)#^Z\^D>cDE?@1>E,8FgQBEUC_FZ?
&,LG-E\JaNg=#_/d:fgXfd4O&7?;A46#T@8gI@?gaX@T)G0YEN^T?;\0BB]L10<,
-Ca@-1&f]5bK2NLY7@03#3\B(FCNVGEI=A=95\dL-4]7F+68@\1YcNcePIPK+IW/
K15_9RJfFgH;fFX+Yg&RS-RH]P8E5OU]RNg)HXV+E7]:#+F[2I=SZ=G?QgBI7.^g
U7YGA+eC-G3W[0Ef8H#RJbL)[S5K#[9.EU\4B5M^C,@A8g5T1Q?AG#P03\Fed5PR
>Xa<)73^QJ=_4D>P<(IW0K\T3PE=gg#2MX3;JA:I/PR22dV/CXOFR-(aH6KJ@>bQ
a=^;WY[9.@^EZe&2DPMX9ZYY)UNFWf/O\D[AMbF()+#[=::dTY6JTC-U(9\OGAe;
>^Mf:_c&>1f:1&BbB-KDF[BAg;NZ/G9\(,&+:Z<c?X><+UH[WZe[_f^E-M#1gA7a
L80(MHBM77DSfUT_J4,6DG;M@V,g]?CJcHRI,C3VXA6f,Jf7VX[=WY?.I1bVF]>B
?TU7Z&c9b/QBg&S<Q9>YHKK6OV#0AS5f([J/E5\K>/@Y762G#;LV[O)b@_4R:19N
0-F;Td:-3IIHG-3Aa>b.Za:?8#J[ODH2U9[<N-89VHbAXAM4+f?0_EGY_@H-AB]a
JHgDg^cEff4>GO-7_?C::/KDe>OBgYIGA5d-\F?Z,@/)E<RN-BM]X;(7I+/93IX#
2_[fLMcg.HLf32=)_;dP4[T#_Y2Y;S;WQ^LMRa6GdcU,,;[T?1d>XVY8<ePS?#HL
SN&YR2[L[5gW]ZP&>1_X5>@@A;^/T14V47F84C)41ZdX0S519<2Y#M>WD)-J5McV
WY-EW\5Xf+g@)GF##:f,TY326d8H??;/AJ:^(]6S2VJRU?2TELXCK90JZNCO&@V_
fcRaaD)bXV#)O1=:gPdW.UG+3@DIG57=f.7c0C<)Kb/DLOQ:(-_>e&=ZLUB;[]MZ
HTT@IE[[P?>geZHYPD<PST/3gUCbB<,5=@f_N991(^RPHeW.IT03RAV&4_LdF2f]
/Z)2-2C3&CBH^8Z.)UZ;CT18&=H7RHH3CY2/5F.)MD-_Z5PdSCeJ[b7X.eY8@(UR
GPc#M;1[0f[^G&.#MH<(Z&;-^[M(:_:=R@-\^FR?Egd1EcHZP3GfVX?0aI\(d:O^
H.R4UX-a8TJWdI\f3>^L#@.H9bK(QZ(:;\Y_a5#&>1B;,;,8W--^N4CEI?^fcR4\
T]0.]9\TFbePf+0-81ceD:TJ+cJZ:[YPR+M4:42^)dS(gB\d(NgYe[f-_Z6Q5bX&
6#C)dbPKeN>e(Nd,KF&[8.Y@NTg6T,,E8_0RRWQ/XXa,_/W?:gLNS_bB[5f&9N+J
,IC[L)d3F=XLGb:LDgA(T]4GeXcOH];V4.4C6d]8UQDGB6<8;A/_CNG:E#PT4IZ7
]d_F&(:SZX\U3gQ#6;Hb+/C(PfVCE&:@RRJ(YN<0_Ieaab[,KS=&J[?VR^a@#&,b
H,<1V;VS17JA6F31_;\(I)1HFL<ZYJZ(CON\0b>_Zb^X7#_--+//+5cGK90IJ[>K
De8GZ1&bX##ZWC:g2,M8DW5MdXJO;6NE0HKFW(/gJ/N.I(9#?NTY5IM7O3T0Y\bW
O7XZ1XGN;[1R:WQ0?;<3]K9b<O-_,ST?Ea)Z5ZWP7<;K5]0\OL;eL<bNfC-L1?@M
D0g?Xf)K,[#<9HM81gL?[b_R6#2M05U>V[<4+&XG]Z2L3[NS]=^[+WBQ05M\XFG(
Ad()+O(6Y,V(TCMEF&])<6Ef4aP[)bBYAG]UEGa@\CZ?FQBH8[-:RM@P59[.\Yd^
VF26g^ge&11@D-A+B,?If\O<XMZF4[1[RX;A/)SR3<O/D/A:+6/]=FXgHCG-f_^9
+URGGYSV()R_L5+75U,bV;Y?)Y.9,J9aQWK;Y4.IP&AMOf<4O<97H62;.dK[Q]6]
RG1.+[BS.\(>9T(_.ORcV@4YIY0F2UHWC+6J3;X1,Te+[NO;@RBGL?8A,?g&75CB
XX2Vfe)[/UB5=f_=.=R\+7;5F2?L-@Fc6/8&I[S,NeUNg-5K>,;6-;#8UV(#P\;<
^8]G6[LOK1-S>Q)?D2DE00,KNAEHd.g>X0S3M:Yd?BK523T4[<\=RQ@/bX[.PQ3#
/+ZH&)4JX6+;KVBS(#PLSS,.I&+)[I82bM,;P@&TGJ:I(9K+W3=IOJY<(._cL3CU
6UY9DbJSTQ<TbX-FJGJ0FbS17LA4D:MTC5M3R#1DVK;#8MX;V[N21Z&S?M:QZ>NX
-gRK-6dG(HPc;U2a=3[GRPR)ST=_E;d#bC4P=]R2X^5,AC&J?L?/4Q+AGaPeD]\M
6VaKHVHS\M)UGP8,gA/Y]_=]fJBEe8UA[b6P&e@&bg<;=[NDVKZJ[29A.6PMI@W\
DGT+D@KIP996&9T_+XB?/D@:7/;3fb#3d7Z/9B=ZAI9T/5KKSC#39[ddJ,-KF-fg
7N)=R;H7Y9IBGC13/?Hgg][J5#\9XPY@+8XY,4c_&4U\Q>^EMgG4_NPWOZCVG<9[
).Ra4NR85Cf@XS9Vc7P?MK#E5e-c57K7Of,.:L7Vc</1M,0Mg<ZgQ[=T^fVXZ9Rb
8M#Y0L,318@5HaJD#1RTYQGJK[Dd[#-cWcU7g)HXJ^+@#,K.H[b=Z,^W2UCZZ.[I
QegfU<+@9W6O/#BXKDS/L0Wf,(9@]3QH#JAaV.>P2U0K1+-.+]0Ne<<&E^gcPACb
_eQ=EJ=U=S-T5E>.#30NCa1J[@3@4;<M5e8S=;,XJW),3(_cH7@4DF.aDX[Q3_A(
G&R687:K#d-FHJGRS6f9Z(>S\2N7E27V?=D>K\+YEgG/0C[]G.^CYa,Yc,c)8VBE
\1Tg#UF+^7>L);3Y^<RO(YGT0X;(dRV>N5NfH8VdEEKBN:E<_PdZd+F@QRd<@J7X
&P^5EE:OOV..c#)>gH_5E+@/(T=N5<2HTCDDfdYVg[?,P_?<&D98S(28LPd=QAN\
NEE7@)M^eJe;c.1f6G5OD<,Re=&O^FSO#UV];+YN,<\.-0YgY_H^RK<7I<c_9UeG
Ff]S,+T<J^RKJcT,DW5G,DgNfVP^S]Tc&5F0A)CAH^RY8H9DD3;9=8b@T8e4K<]>
>\C,+C08.5>dGT&LJ_Fe1Kc,;Y98H3F]UdgO>6>=P1U0GNS:M<Le_HTNP:ZP,[);
f#La:Ze=]>WDJ-9II--.J&U&:@1f.>fUNCHIAaAEd;5=JY>KH3LfV>)@(W9fTf4F
;6<-.E#\5_654;.PH?>^6^f5eE0fM-CV9]X+XZH>.U21cQ/6J6LcF/]RA<0Qed_O
g.2EbcNAX//:]Y+D7<45@N485T7C;5V80CI502^9&LcZHF^aSaL,3d(37-?MbC^9
<^8H8e<fM6FIdM?1g8=@#FK5](YML53FgG)9DT5(^b6Vd<;J5PYTQ90Z^U[G^+QD
EO:D.-?(J8BD3ba2:CJU/::W_W3/NXQKYCP-ZW-1BEV<b2RM[^M#4KJLYO^U<I9Q
cVYMXN-XD<aaN^SFYT.6C]GFS]eG.D_@^UU_VH-+^?YZI(R,FJg^(2#5F6][\S3L
)EM:?&DS87a6S#YV2WUK,5VaT7=CE53+=VM=()A_ZK5VH,IB.IGag+,Hf\[MfJJY
W8X5,3,17:+1R8FDf#fYMZN0B:Q=gKC\RC(7VEHJ(.5==JM5(IOOAD=XegSa_3<P
0OD&L=B2>+5Q0cZJb]0L75FX^>YPIZ?Q;2e8B2BJFZEV)8RSL7-V?fSgBc<@U&]A
d>G9c#c]&<RPJZ<L[04]92eMBbN.S+;^=R\A/HP[4&M6FAGA<+1)_?L4HKc+_28C
WSY>=24\Y,WG/4b,#d?GIQM2Fe@YF_VF9(8b9F01+:aS2KUH_BN0cSeQ5T&6@Y_6
Z^0LNOR+S39=1(E1a.4ZH+X(ggJ\NWG)RIF3]YWZ,^F<CKeBB.;.;NV@P]:)PS7>
SCX>1:\QX]46X5bK,4YKIIa9aT/&<?MB&/KV<R+&F?VYA^H\F2]ORUKCN)JAe<JP
B&]7d2\8IbQ1,.Y_DaIf]CZA@2d_&E#4)D^UC..5G]#3(A:W]d69+Zb1bD[c9b.+
F3,1WA[aWJ;K;])V[fG<\]#BOKQ/B?@B11B6N&EGPIObAVgbD6)Z9-98Fba&J##6
+d@MYYQ6G8<>P;D2J_JA_,31Dae>PE_MK3bL13dOF:B2=+O1)#;OD)E61](.<dOK
A1PP(6a/GFY.US036BKRAQLKQ<<JgedEdG+H)C2(:&BL,.7SHM-8e7EbdVY(,J_1
L5.U7Sb:XMQP:5L:]M&b1Oc5.@XU@VF)UNX>0,IL?68RMD6/H3<U:__)C(5g^APD
eJ80)IbRLe-JRE&L3O);)@Ag6FbgP96e6#KZ84A^7+.g&M8O@24S_[QAGX@F.@S_
UB>BV6:A:^f62K(T3EK7VUIcLEWfGVd:+1LW#ZU8V88CE<98:.<;X>gV[>^4+Y.4
Z]0@VMA1)VXKb=QUS/-1R[@HGLX).&<YeSQM;Xcb(Y=9KX?.\)N/9L)FEN<,04_B
TT4a@M<F;-X.-3,.PL:1adN.T?T.5VSfe>dgR&YVc8e4LV8C;;Q[F1UB^B^4P>[N
\O8+H=SQ\=/2K)gON+TX3@C>g3COXf/RR/CcX1FUfbbA&.F52N\-P6)g.)4a(-Fb
3I@PNI)MfbD>V?^<[,?AKN:SGVRP(XKeOYbA.38E;-6GYf0<:@<:PUZ900#VS@V6
W7Q-X/<<W3Y&@MZA1aD^I2XQK#(CO][K75XI;GN(F\3\P3Q1ZF9D?9ZUG01,LN>&
RMIc+.+FOA/]<FUe].A7E^GcO;0c=9Fff7/#<W[M7Z>d_FT8<><32DUZeHU0U4>[
6;8d-J(]Q(OaWQ&U(#E,eWMH1-WEXM1cM5)LTAMKLP?L>9^CWb4+XL7TCR1:]X3N
Bf6b9W5E[#]e/gRKXNF2&4WG;BCXCB^D:?:\Bc7I<&aY<1=TO8.-gW6FQB\+/KAO
?f2ZeC@3?K,F@B=@Ef5,[VA59,3CKg8d2>)+a^:JHdB#6@M1Zbf-gKP5_R?-V3BA
UEFV&CS/?:G1_6L.Z[+/I::b2Ug3/M87&FCNG32_1UTMH&(N94?YaN2KROMS4S7_
XI+6Q55^BJ#(^ec@Mb,AIE,I;15K90B,KBU<>IB1TK@fL]&Ab]/F.7Q0\[RJ7[A:
-T4&bQ&B8QQ4Y=-1(NEcO[R=XH\B1@;6=U_QQEQaXX10/2X=cXSA>K_855bb\6KQ
a1ZA5O0AFd#J<#L(gPMc;DPKbX2+gI-_OW3<=>+(AR,4g@a4aVO8RCAR\d+0Hb+R
8WTM6gX(;_TUT^8.60/:HKHJT^F_beWJSe2JVd0M]e7-a)=,Lb[-LbYaTdc_60&^
[fBRM8dbD0[TYF(FJ-EZcAX;C0NacX/KVWH9?Ne=]5R/BCV)4&.TTfS\4+1)KHOO
2D(b[KN?eY9dG<HTYRcdJ@0_?RbJ@ZK;d8(-=@WZ;T:GKN=>aJ0;AD?T>UD/(Q/5
\.LY8,a&2&A(U/2/a::D7WU@@J4fZ09WBIB^/=A]48;(5P6.bE6?[XOHY@/J#)IP
0XKdD\28^NSe=&;I[18EKQM2MOdH#M[+PbJS1:\b]4]-IB>)E;DZe)C^_A>BPX(d
cCU;F,?UCAcHFH,2:6RB6G\5[KCKO[J/O:ce,f:;XUTf6d;@ZD8#:P1&+&TLGT3E
M3]DC-[gXVG:_2G0B[K<e6VS)Z+ILK#^A,B+fHUgBM&;C;@H=@e\9H[VCZ/BAfC/
\0gPP=OPeWP<MC/a[f/6][;d0#5V^()(:+UQW:4UeEWOeD?7IPKaORC\AO_U[f5A
aF6JYXXMN5UJD.;fB@=MLC/6d+T&WK[;ZDdHFB?1\F#.U&JCAKZ<2;#,[E9-3I>b
Z_D[E[L&VO8]e/2SQ/NU^2-b9F>QZOScG,U0X?)ZS&KUY;G:GZ,IJC>JcaV701L9
bN.L=cZA1;MVN)b-2R]=F[+c:4Z5C3O&.[S^dJ^Oa>11:If)^BS8A8OOBeQEGMUA
\Ig@DET4f>0ZZG^cY2G7U>(14M.A885SKIE+HC?@VDa=ZcG3efe:6/CWBe:-)Mc3
-;.gJ3C9/0Q?)RE?>/9PH2+@>;V7a7<._cBd;2X>BK\(<NI+P/d?Rd_f606f&58d
KRa?\2@g@AB<CZ\ZfgR5N8;D<NIO3)[6K^FUD&#8_Z:^J[J]fZ^\Z3;KWOLd86NO
9;BF3T>QEVPA_@3U?bO2G@<\NE=a^]],+0Z+CEK1\,X7_SCW,D@g8bP93f_c8-Y=
;?UN:)WOVS&AW<]X;^BUDG6K7WQb<,MYgR&_-?1V-XNB-LXV8[7-D:TMcdA[H0&c
RO;OVXA:Y8)>.])TF33V4C109YV&OHPeT_/cdUdF_fN8D377P?Q+ZfORbD8aZ2dN
AE+ZRE6ZZe[TT[JU85[E(.<&)ZV^=4,Ic.D-@eED&C(GB:3\=<:IbB/2U;<6JT4b
X@[NS-MR@FI9\A--@b?[2<,MbWH4]JP=_23SFOUR4>3H1>^@Ag.),H3aIceC[EL#
fH]b=8PdHE-9IJ6U)@\GM0RJ30GAP,d^3@[TUY5LXaSZaTN8VCg9_[Df71MJF87/
(HYcR:CM/@[@I.=JN>.WHZ&_a9@>IQ7,Sc//(,.TFg13I(P.f;?7=K?T\1VbAQ)H
,1bY#3J9L5C,.dVRG5E0^GPbWG(ZR(9&Sc4^ZUC:-A\EH[8;CJe6,SC]O]--VYQW
/AQ<Z#^26.dL+36YPBG6bLOQ-(7>,^/GJFb]^B7I(YOVM0LJ<);I@=YXLO-?7)fb
^Z-[FMT.0:ZNgWFA4/N0K#9DWO8;PQ&V5Zd^F[52+U7@#c_ZW-K\0Yc^BU+:[J<F
-]FIddVYMW)Y;.0TXQ3I5&&M0._0VB-[NT4H\dZbNQ5^eDWF/B=CJ#>,A&VQ;e]]
M(<)HH?7X9c3>OW.IF0(P.BM61-;#NLaYa?;g1TR[9H]FM1&D8Q;\d8gIg:S6W?8
L=B:e&9dXd.8gJH_[f^?#fL=NAH=fX6#7N+@d)880;>-_QCSGc5Y3]LVYAPG1-Ib
RE-gdaBL?<0WPQ+2^^:b_c#@a/P\UgX0g4TC3LK_D\TAHB8WOG<BR4#W-/ZeDeQb
>K972_AS,?aV02;]&3GV2<IG6QXGbI34&a8.d1L<E]^7Y5NN([MFR1T>-C8:7U\T
O+@,40@216ceYWN529BH4cB2X+?e]:d\Xe8@T_654F\8)a_J7-)[VA^1JJa_A25/
D302GO<ZJ:VHUUGeI2H+aK.+:&?D+7(0X;ATUA>CffN9,aNJ5([WM7a,M)[a_UMf
26D\+A/P-31G/FB-4AJ<R7[fM13C>6_FT6(WBI=X4c)HD@2WC;G>=6SZdU.N/YIb
T?3IB0NOC=dLfN<WQ\+^&M1]=8@8EZ1FR\FA)R.KKY?M;=@@d8;/TRb.W0\GQ2K#
;I+S8;MC+3Xb&>4cULR12^;bH<P/I+>M7XE&APQ^E)\d/\TA:VP8aE+9ge/<e/1b
+X;)QLMK>^[F54[S+]D]U,WTa=M:aS^.4@0@(U<M_?f0Jd</>UGgRVI42>HeRRP0
[,^3E&<\04PL+QcD[c_CLa6FV-]S.=&0ZXQ@[ZD)KV2LDN<WV9W9ac(aO>BTAUbJ
2a&ZAOG.FbR#@^IGQ8_L>&/DTBI]WU[>AE14L[]JA:51OUCY/PNTDT:g8(B^I_]/
Z9O]c@8_;G[,e?Z,AE?&9.P^<Q;69]_I=MISF=IS32]IJL=E>340dg4,Be-I8-aK
C5N5M;\HLa]bc=8,-d^PX^QSd6\H#/:LWOLHD7B?);e=Sd&ZdK,Q.:;a7@>&GBQd
H&XQMN_ZZ\PEZ87A[\H_57.[fTf\TEGY950]/)?UTQ.FJ7TWMIVe)b<,Y>^^9f.V
K>-IOCdQF@MVWF5CdZf:aY+:_EdbJaI<MKMWV&X#MJ@a/a0aH[ZFI[XKe4>XMd]\
F:\:3T:W9F=PUD>8g4>=FaL6/??YY-FP>_/QWDGNZGf8,SYX>5D[#7_6>GOPAH^+
UF6de-/^83VN8Z+2V(TaKYH_IaD46HC\a=;5S(;#52[JS&7WVHTW4SBG^#>7RPC#
SU:eFM=Q;;3RB&b>2]M2gM(cUK-N#\6^Qc[[X[W-C@3_TT7,?.d])L\TX=eQb]W;
PGV?A0^F01?]?1,FF[g>-IedL5;TXXJbSB&B)_GV?TNbMfacbB+P\;Qg&XdJ=:^.
6&J-[;/Dg[LHNM:MHO.DbV<OA\g3NSPD/L:eC)V8(#PYYVPagT+8BfEH8PcJWH5G
gQeB+,^FMaZSgbIT,/\S69XIaNd,9L\901aKI\J;TQEMO/;bI:e@0LQPE.:gK9?\
W+_B1)g\EFMPd9^DT\RDU:6Kdc,Ag#;=TSHFAXG<9DV3E6\\HHZZaPXQCQeEAGD0
Cf.IUSD^+8XPFV.399b,g^(]./&YPH(0^=eFZ[I+G#AKJ@;1B\3Y+?;[<I=&dcIG
;B+L?,GRdY(d-TbfbU3YZWb<A=0\Z#9MF@_=3HK;Jb;AF89=7OJ?MVC]aOYL9&_D
BJTMg/6UeS;XbK<cRb8EVM4NH[8N1-#T5IZA#7<\H6=I]MSO2HR=\3[c;56Pf3/W
ARNWE5+-6/&32J00N7dI(46^^3].@\@7V5_T]6CF-X0\I5GYBLT;(#e5f5aR6D4M
d;W8b5XSe?I[+:4fJ7dUbIQL^5MKPF=S&J&[Rcb>/0<7;W=9(=8gQ@e/8C4f2,U.
[[.eTM723AY3>b_WT_5_(3IW,1T>IC-;G+(AP>cg]D17LN<7:b#?<+_d+BE]0T&+
9WY,7@T_S-2MU7,gFT.b>CJTcP4dAb8@#)?@9L6\1)9E;fU>_3-G>c-LRJ5<Zc:;
6fd--g0S9V4LM,16SWT#O1\ZaM5=#eS2eg\04eIUH^YW]8Q-@,3WRON=B1KA07T.
(GRC_0^0&XRWdL#(X2=UW2^Gd8LEZB<A(Q^8FFY=^Q_.2,:e<RN2G2E0OK_F4_P6
WUe8FOXUAPYMaE:aO+IF6DLD/.QXH-SN@&;.K+Hf8#5OF-+ga[+_>7S]=dBX[X.a
NWOaM:BY:b[4;VOJ1;2382U7EEP-1K@CL.L+=<Y7S\6_PZF7_DL&d(C_Y^(,a8a.
)H#)Yd#A3XTJa,Q>_BLcV.NWWc[B:AV1\e.dF2Q;e>3E=MVc1<>9e6[)3TRJLU3?
\0@M5/S2NY7Z99.CQ^IJDX1&YQ8;?;9D(P0a&=g.^TYf,HJ]Uf<2FCV<#>7V,\:D
ER?edOIAA#dGLAf)28Pg8==Q1G7FDeTEXcV1ReAHg-]6RX^UQEX=TT_R].-.dGB\
eN:]PeeFYB2ZALEW[5+Z]=[1QR_MJ-IO>-8FH(c^W-\YT/E;5&\->_0J[=d[eH7L
d3[af<dN3EW;QX>RgS9WdLV\0_O+N6&-08c;ZNQfP0MNU.[UD>;&5=G(8ZG8_C(9
.DGPF)?(CCP4#_PRPO/:MUJeQ5QGb_RIaLML3G-aDO?,9UcdBVY_J96Ea)KB2=aa
4X&?+<caDF.-DGBIBDFV.\&>?Y1S#R1Q>&2?]V>7\eB>M[g3JM@K]cOGb=M:4<R&
aHCY09IY>;gAIcSQE@C]K9XO;Pb@-d>dX@Z2&./3,6DV\BAZ>R58_LYA[1<a9;]b
R?^YR>X0BVT6(+X)TZOb.JU,]^@MMR@\b;)3(U>+S+\6/>D_d>=Z:)IFQ+4#c.?D
0dYc15^]^gPS)2E1E-;&M9<8D?c66@.Y)@C[^&[UM3F=?:Y>SJF2,c5?2FNbUG0f
eJZFdVa7/6P+]KWQ=<KW6>cbY#XNG+gO6D<+P(#H6#=SNYZ?S,2YfLYXG@Sg;ZD3
JY,H:S]/:.>TU^@T:X?4U&c;EYO6[EB)(+C9,V3I.AP(<?5Q^M:<=g1eQPN)efg4
G@LGUO<Wb3e:U2:K<_;IH,4A0P44PQJ,E:70C8U770_PBNFc7:-g.?Y5S[T@RW3+
3>JVD@Y7RN;Q\27b#4B9-];_Jec=7P=Z=FLFF.,GHMDIa-PRVCg5c[Y@_Vca\[13
cNF#?A99[^=<661H1\fDR,&/]0<C/XBBJ30<&Q_C6=QRV;3=NX.2+?Y;V7K\U=aU
/f)YL</E\7Xb;4/gBBB-;.\;O9?_R0),IZbe:^1W=dc=EFQd&>Q./2(FK_Gg.U<U
H;8#10HS\&7G?=332@1I;AaR(9YWdCA@a24#Z9VXa&Z.4>^.+bFY0#ePS^78MD^L
_:5<8&4(2#764Lb(@<138>>IR-.EKQ?.3-8@gJSG]b&TCED\(#:N35b4URW+-&/R
3#-(B^@^L5H-#@RXHc-<aF<c_DH9(VNEU2YLC38d.@8.@\,76X+D_F)S?d6JIR?^
IJU^S>+NN\@CBQ(W/U-cG^fH5C8+HAg<E8173SWXIeMM_bU.Vb#f).:VZ=K1V<;H
81)Z>3A_GK,U8/#3]1[)\Q[ZI9b?M)=B;E>SH1YIX]CAC0I1U<bX/.?DN-[-R9Z^
Wa0ZM:./WbZG_.&&>4b#SXY2CP0O(#UbO=I\_a^H4&>/L8DF@+b1O8F@/_5&-@6F
WUH:G(U+_G58O_W#3c/<[K,e#PL=XKP=c^Ne\46c7072TJIaXfS.P7;G3@DA9&(5
&?X?::c8#4W;XJRV>.PW?N-.f[\UU5B3<agX;FN=TR8;W5P(EPG.CBDU>SSL<#7L
+XE,^,(AfaK6gFG=,cgQ[Nf/9_@a+@?B;+ZW/D?d2?)RHd39-RLXaZ_;_QYZWIV>
U\LCHX4SVHTTdR&)TNd][[6=Ng6-CM_YTe9>/;.:HbC_B)_La51\=VFV-bbW-YbZ
@N[2/A[gAe-e)9JOK\G?8P?J<5Bb-]TR.X\Y)?-Xd,^[-^,51e[YA@N0XJKdb=(X
GZ:;U6???:R,a3YB7MGD<E;fO@TWcfS,B(NW?+8I5=,K]XeAPYZ,RGQQWF;B_86@
\0b9[56DEGJ_:.O@?0P@.>=&+1;Sg_;O62.-S\M>Ja&@J4Ta9b-SDX+)dg;T)3W7
9a0J/NHYVSP-4Q.[&3@XHdJ_4d:2ZT>(<7gMW_B,+/De;M\[T?NLRcXQc0gNQCMR
ZI]YZLGF\9(b?d_@<YV7^4@/c]_4e1&H]O+R?UYZ>b1Se./e[_@/BM_>_XHKf(I=
4-I?L[Cg=#.1@6.6+AgQ<;0H3P#_]WB@._3M.P@?RI/(4C:<#SZ-PW-:Qg_\M6SG
J[2BL@YWG[0>J.73M[aCMT7CLO#dK9QG;WYa)7:)8e5^-DHH.J;Z0.BW^XE@E_.#
=9eG#X)4C#bU.^45Tf&DEb4AA__VFMY,ZH:^Oa18[H?5ELeQB(4S]96D6SWIR>]]
PT\O9E4-6<e\e@3N<)JPA]X:31^NQb:YQG=(H,LX:KG_3+-c,#g2BRD+77(]5WN;
DY)Vg#M;/+ceNQ_9^^]6Nd0fQE\9,\FN#T/,GU[/8Gc\H+GC[8QWdXO4O#\.[O+U
3=4+=Ld7/0Ta\^f3#XET#5N>SYT;g332Pb&fH63AS&A?-)GS7/F2FMPH7V3-Q4@9
<P8L1OD:Pa]JRJWF:(2>=DI_Y]\X+NRVG]85bIebg(IZ7N3R&/aa7IT1#=6Y0ScD
Z[\W)76-@b.bN-.J-8W[K_K8#I[ca<.b)#Z;T\fO?EV3+:c@@RbFXL-gWXcMH6eS
]K.L9c4Y=O#5/GE_aEX8>4^JF/gL7PC^)fL\C@G(BPDSJfM#UVd8Jd@D,&[4Q1Xd
@PC:QP)T[^BYI=N[ZM)?NP:#9K&>I0/@Z^YH:SGX8Od^E?LAD/+31<Kgd=KNccHS
:QG#9aLHHBYHS>\2]P?Ee:=34G))Se4:I9JDQZM.F<g(M,ebF/YEbJHHf<I)#HTe
XO6a[F106^>34Q+@3E-Q^3d5D6DDG8V#STAS.@/RagVe6(KG05N?g03N-EM\;QWI
R4I6.9S96XgB>1bWb:NJZ<WE9VH>UVW--?[]GNT<IG)8N)-.)_BXPJ_+P:)F&]4/
Dg6PS4c@G2<d.-(BdOJE(/]J[c:XH;&:<4XG@D)(9JSWPIVWXHJV:X/J3CEPL6:A
C,d_ARV=39cYFeH:D@90;Ze_MZ3V#<30Tf02b0YG3DJQe:2?F[DM&9fJQ#94QX;L
U>Qc1ZO85?KK,:c9\L;M(gCU];7fb]4M\==Af&IHVZE]O5V+:)+2//8CV#_?IB9K
U/Of)gZCX7JYST::1IdBM-U&75FRUAW2=R/QaA3Na-OJf@2bQbSCF#(/(^8?HXW#
[_56/aW0/7YKefG7O5>CC5Q_#+XW^c/ZaKUVXL\IXTODd3(cg2,7[gG+6b\_dVgR
<C9,MRL8\-(d,H6)ENc8/4(^=a[OM&]]=X+(.Y82c\cAE?Ga>dbQL/f3Z/df\58_
N5^Y8QWKJ&F+/\.Ebag=H?29TQ2P+_>ZH0&(Kf4Y?]K_WR5UeLQfffId?0FP][BH
Z7O<5CI2(V=(@YcZS+1DGb?ME(a@&O/?eFW475.)FeP_3:g=6[,E_:dW^#a-^FWG
2W+g>M,aR;Z.LeF[]A/b-NBJK;A;Q04/X.O/@A=@W;?X3R#F#f39cgK>f-0;?:^7
&.1SEJP\\JJ^)L@+E]YQN6I.)UR9WWT4ZGcS;K\\dU<WC4O[^4?X_D/8GQB[CCdS
CA+>^2_#K:3/ZTQ+_@HNP6MB9HM[eKe5@<@XKF^Y7_@IP[::<?&=GO1OTFI4:aE_
[^Q:PODPRKEIOcHD]TB^DJ#FS,agK)e>CeLS/CbK=V)OGEP##UFXF+P^L;O+a,#d
.D)EB&O=8fM@J]D#A/<OGSBLaEC.UOZC53.1[e;Ad4MRP[G>MG(^PG&QHM.@9cN@
D6XE>H,5\;W4W9D]OSJ1-5<D:30eW8JZDA7CffB1@]6/0:#_Me@b<203RE+G6OC_
AWff1bV1I32dLY<8S,E_W1c6H#M9aIXaE>_B@04bZJ1F3>GXed?R2Y29SK_Q\JH;
F20RWI?HeJ0c.>G_gF1e7))\#2I)OCe=\ZGI^VVa4Xbc72XY()I8V\<B74Q3e7^Z
I<#L;HU6Z<:U7SK7d[c4;D7aFW,P6JdUFOTb>b//(f;33cO3JHK1RY1GVK/[9aD8
[\?SZ>4L+9LdBUM6O:VRZ\9()-E1.M3[@W3;A3&(?.)2BWLPFK-:6\V,/XcOE\d8
5aT.D628263L-]56\T[I#F@PbIWcV<RW2e1<I>IBTG:7UbREDT:_+UB@EdQL<7#0
3bYLL>bJUbJ6W#)MJ>,@dPG9IO221FKK(&JN3&FUFUCW)e\D][VR[BZZ7cN+R#])
0g^O?+[>-K7W1FI1];g<SaBZLXcEM\<(bg8]CK-g/2EM&fb.LO=0Yd8J8>Jg+:b@
S^6B6SG9FM/)?]:+=PFF@ac]U8CXU41.X.be)EG,8<AYBcC;;6K+D4]1].E/f9eT
JNge\7(17&X,+BK+(96P7+,JHV:.XV@g@BbIH0NZWXda+U+93^1]_G/b3d)OfaI&
^Wb_bU6C@EA^/3;1F?TG^fA[X61#G\5Y,?TF3>MWcT@b^Y3g0/YTc1-OaEbf6/_?
aCK]4T(agW[]/9QA0EY@+L6ST.=A1W/B\FL[(-3WRXK,96)NXAa.abGd.\&F;#Y8
-;P9-fgc2baS@575C7Y(_gC8?61Z+#R^[#V.?gBBKS0Vc(B/ZXH]+XR5NEGHY?eb
@7?BbV9R]/N=]95a]F,PMIN/N?,\FZf1Z<EYUA6_K_4:b-1<UAZDP88^0d?(4bSN
bHXN_H#--0I6E3L?Y,A/:5)74Oa)DG/T@dC\b=K&\d3LV,^UcZD]4HM=2EYc9Gg@
EcNU2-H;ET)QY].0/>OMLBPOc3_1QZ(FX7#]_2bAcb6&La147CfL&cQEPTaP+V#T
2J1KfQ<N6E/WSY>-SPG5RVFdL]FdTKL/5ab3PZ9NeYS8b&.-58NffBZC/D[+M]BR
4T;.#.F,d.1Yf-U0LPY\LC77;_,,ICB+.J7:<C[=3e84dG)8aIBB]DE)[7dY_QaK
e^#YB?^8<97a3SJaF^FJ6ID+SSaY1dWXD7JX.1K#/E[08;#d_gG&f1<EJKY#)?>[
@V_M7NaB3]>>R0:I=d1ZfT-AV>X5@E.LO7K?_f5HUL2D^G/8>DW5,g#4)QV]<^@9
JJ)R#Z/&;Y+fd?R-#;<.)WSVS3&@CMGS_0f]L@I7ARWXK#FWB\G<=MYQU?D/CK[g
WbP(O.AW278g8L\^4[(5g#J36)3b#<R6_AEVA9SRJSKBcS@N+QUI\MF9LR]8b:FT
&[9e51M+D)2HfGf:+/eYE?KddB1BaY3>LJ:-B/Q&.+;cTYb;2^GWL7YQBd+WI-PG
VAdX2M0JEIS-;=T@PI:SOQ1T]YQQGMd89\UPUgRXR,8P]FMH?;?AB[\N(-LJgcL&
.O(JN-8<9UJZO.X<@PZ^&V:F9EE.L(3UF4Ld6JYT9Ye0KKdcDGG;TL25[V,.<b]d
gPfL&XH(=3=9d_&5,D?G]g<TJ/3Q_>TP89Q?BcCH_b3cZY\UL@ZQ()Ud)e^9-XWL
+#:D1-3@7Y\DaO>ZY,HSHV2fEO7^7X\@@_3&.8>TbPIT,V)4YOH=@IUOMgYHeVeI
\BGS<5_;53\#Z)S4D=1-dF=&/BTG6UL,V1E#?f3PG=B8JPYbgE2aa1C9cOEX=;/W
e(X7d\-;5g;FaH0P0[JZEQ&C82b719c#Q),@X[T=8becI;OXbd^ZBc6IdNFTP6?@
G+AT5Y01:@Y,JbO2I5/GYJL_?31/)HUAaOZ_E(RI9NI4C0H<EU0HR&Jf[L#S-/cV
B.PAW0&bNU=Bd@EaCKb9R4(AN9,_@4N]Z@<>:,#7ZF.4P=DGXZZH6-&cX4XOJ3VG
]6G2X3N(9bc=OT6/MP)B:CT4]Ef8]\f7b>^@WOK2Z<Lf=#SGM9XO7&DC[Y]543^0
PYOb38KV\S#ZAQ.A&fF(bgb#A:7<0O;[HJ5@PG4eHZ>K7V>CIJ49=GVDYK3&P7C]
.eOZ47W6GgTM)QEPfJ+M0&VC#5\&9P@@K708LA26;2fcCJQ1&J^XY.TEPQgE.)7O
S8CG;476W6,@#NMT:3I\::65L0:a6a=<.g7ZJe50Uf@#cFEIZFVO_0WT8Q+dEHJM
]Za:9&,POd0Hb]KJ2U[g;[,^b7OIEFO/;LYGV,K5Z2LIcU93A9Y#7PZG(RP2dNR?
CL>Q_@4Ec;H#9D#Q,<&IIVT6,f=6c.bNfD8FI.&5V/R^Gg@cPLDgbU1ANfRR4E=Y
H^d?\(&U0J4fa7B#GFI?A.0:,eMS<K2Je484AT6d9#-_4W.Ef;NA<6>4-NcYM4f:
GOUGMJ._SBcV>8Jg0Y-OGESGcT88FE^DD:7]IP?HC+cfIBUK2WLHJ0/H8T&[I/HW
A_(U,_NT.g-)Od8Q1BOfF\--)?C.:dTW(Z=#=LdH4Fe7^JA6,a6@B.[@a-3944ZR
ObFW:f8.997]=>>JM5DVfS.IMeW:9K5>=_&8&(/>=PS[;_Pe]FLg?:dS>gd1#RXV
=bZ^/8WNER8VO+RJ32^]?#2VO0(.>G7\HJ;2QO#2Xc58)^Y)CXIRGf67ge<A8,VF
ANg_+TgfXLa^.QOUcT:\cfTcaXb).cN[N2M&+IHRYVCW:T(RgO)M#d;&(4Wg_3(J
5RJM3513V^N.:M;ACVF=241MY>bO+A);J77Fg>UD>HGZCgH?GKWF-=KO5^0]C@Ea
aRN].+U0M6AFa4M3Y;=U_;^c:e#c_GJH8JR6\\KP7[(Q&bG^-6c7M1@-6&\)\Q6J
\d:U&5_\b<KX?gI[W;gbY7.,O7A-/&DRX2TVLW[P_cL_;)HXa]a@=_]JSM2R;O]-
30@9(e;W:&U]J[E)XV:?G/AT21F[S-N]XCafbT?7GUeXXA3P)-=@.4^-,^dA.fb+
KT_^#Y60=TVQF2Pb.?(5ecS1(R&4XLfHJO[:I@]=1TW5.bRHTS7BO699HL.);FdL
Bf)JY?3P\?/S]H&(OK;2&9^;CP@\d+AafXQ-305NVPS7=@CVQVO3[6(WX4DHW\fG
34X5Jb?4#\#I743H>)g/B4#<#AF@1Q.KdXU+CF,>-ZSa^S:;Jf;(,#K-/[=-8(>d
=0JN),I(42]gITOd5e^7:AWI\/3IUJ&/Y1RB\ZTSV]Q7KME_UdRWfW23,1b&B2?e
3Q4Y75_X:M&O\=E(0DI_fgebD618X,(dD)O7-O1=AV]BL;XR+;F,V_gQ2V2BUPAX
Q9(8=&g:Ge\+XW7(ce&8NddZ7VGe=B3,Ca::8DX27C4B;SR@/O3gVU]DTG:?O4:2
P-XC@N,fMV=\T@4QdXaTH<L,L->CS/C2?V5QXJY1;f@8&2e9PP2bF:I^(B<47G]^
e2G3,;Gb:1&XM_>c7T8:;f?FO51/b>)_N:>fJT5ffJFb2d=[2(F45;e4)c+TEALU
1fD4(W\fN^\SHfBaM=DVP:XDQFULd4c#FV1]7-7W7He5R#2N@NQJ0@&J>VE<GI2)
&UAaU2\9RX[V6)=eOVR.UU-7+R+SeFLR-Y_0GbN>5[Bd@84[4f)&XN5cg,B58Y#<
F1QcMDV#ZP]UfXEZd?eb&V=/X^2:WAP_UU,D.fc2AZI[.D.0ZN1)/bN,2\OV]//+
bWKd^<(^#0_Q^0.;D-99#M.)8/7NEH#ge23OVQ;I35+3(ZC6QI/A;BW-3@-Y7JaP
)gLDa:,gP\9a@_eHHP3gE-P6)Sd9IPX;B[_9Z^MYO7GLdMOV4<\T^4aHd]Y?;IQf
c1OacM5Mf9MTg5c()M?W=bU<,Z&OcV0Db[_5fC5L#I=0Xe(B?4^P4)IC#5J.)6,4
\Q7Q5F^[QKOIX455XKeTg=6#&=UOQMC,E/1[C,bPg3/[e4Z&gE<D)#+P^GJ3N4d]
ZY+Yd12H.3c4(#f;Y7=644(258]5N/36Uc7<T6+].0.2_Ae&bVV=dD-O+H+OT#Q9
R]/+N7[F]V,3G>H0T.Pd@QE#a^<NBR_7a6:^WA06-Q&fO3VTP3O@9VAEI#+BW,I9
SSVMA2C]3/UYd_]]2_a-La#4;X3[+PD?a+H^5LAH7,Xc5d#1:He2P2Q:,QJN8JVV
a[SSJNX/1+LF\3YLAOL,23HFYWL3e?cd<eM8gNg=QdAe\0KOZg//JN2UIe50S+bH
<;C>4I+809gS1)3OA,X,RD[eNZfZaBWFX8U:48)R<T6<cAYRg8cU@F9?d,@L^QB4
^R-J__E_,9gV.DIO(Z(@,/a1A(5W,:):07B)^ec^24E_G8>JM0-\.GR;)<LM&fcP
ZY3QdW@(SW=Ab,Q7RWV,,E<XaLIWAaHHcXZMH1,b]07aE.(<_38e(W2Nb/3&K#?W
[cf.J+)R5C_QO>B//)OE)ISaLa-3QZ;?bgT+@3-_D]Xg9Q/0]Gd)-Sd83B6]ZK-d
3:fTB\ZebEXdWZ>@:.A/L&V=EeFZJ6#8/+74b)SI;YI\9Xd#ab?f&cY-)VP>Rd9:
7:/LCd.+PR_R0J&=2]6T:3e7I#Ug09C&_2_/?@9aAOX-aZC>(3JIUXJ7<KM/(_N>
#OIIJ)(3HI>37Yfc?g9O9FGd0_<0MI7A5;>Z[-TNWO0c95A)F2,,W[SV=Kf^30IY
.\+6^;5cN6]>gII+c,(:GG,cQ[AI>_6XYE&D4-dYZA:dgV#:U3<d7H;WTN)c1K]1
>;?-M.SW?U.L4@H-&,?C&A\1?E<QOQ^:U>8+UXM,)-RZ<;T6<a6V@K1784F\7?c[
5W^+J5#A>+=FR8I<I.4Gg;T:IP.^,6I+4Y-2PX9\Y@eV9MCc/M<^f/3O;56QLI#S
dE<5>>=6b48I_Id&(-\S;X(dOFUJZQ<=28f9EXB+;4_(X@gQMM/JLO)aY&ID+-;1
b_J+#\,N=S>0FPV[@\]J=#:bYO2--Y?/PRS?(Fb^?<P=cLF5@We)(1;((T2A5e1+
4g+IC+,FORDD5O6<Se6.PUUc0#ISU/Zf&&df2Fe5=MMc5IN2N]GJI@/O@KfA_[5J
-B:(&EAe8(+eJHN7ZY0Qf(_EO?Xb+QcU9Ea481&EMKF4->:;891X5ea^:KXLW+@@
;1_Z3=Y5C:@&-S-U6KHAL:C;1VU_GGO;MSGF=8E@^8FOL)9GV/=g,M_VC<d,COZ0
WNJZc3__DMaCf\DaCc9O[ANZ2DQVMH/C#14^dH..Z6da1/.O8a+,=M+QF?Ib^S?>
:,3+7?eUE6:1.Se.SLU5KAY3O?G&bN)LPJ52&[[&?S81+&6d@bVGC#\JE#4(e-M4
MbHY9Mg22F=Q91-/A3)84I.68>EFJ6PPQH\#C@A[Hcfc2>]3Y.F_gQOQb-/.&X(e
@9^ZU@fO^YZ,;f#QVSKN.AV#]7H(Afc/)c-A/=TITF=.b2]cOd_/Xa<c-04/@bI_
1>a>3_99;A=c9,/P@W7d?9XV@>)I&FQ-Y5)R;X<SOIA(4-,gW_L4S^TG/.8E5]4I
aYXJY<9Z>F7Z:DQ:#5_)=@Rf+L72cg8dTH6bcW,^]L/Z-:BJYFS=&F__+PF((Z\9
IJ<U=Oe1?KdOT:bS3H<fGC?>MBUHd08OXY92U6IOaAaF-&cR>M8_DVE/_WY0CN9M
SZ>a@:X-WQ5\e2-VW6K=.+:3e>RO:84eUYWX+KXOK_WHUBLEPb//H,:?Y,(9S\JE
#8&QG,B&C(7YL&gAQdfQdU;A.1R<1gdN<g7\V-.KT.+OMG63F]BD)eF&7E?77GK-
0>4S</I/BMVO:E)FDFf-Y_UM7:Z<^F>gS0Q3GD(=4KI_.^fV,#-NCZf2<0?YXb\W
DBbaQYf>A:__JdXCBE,)^AdP?MC8#Y]]bcAf?I@4.0-a:M#^]\\75A_3^]2I7)\(
H;01D&OAUE5?A,NC.4J?@aUbG-)6AI.LPJEUX6A77IHAQY@UT=9J23LDZWW@&[Pd
?W&]KS.7N5+5a,_K9&#1K7,R_d,:2bcUAEaN]ZJTNH33A:S\,g1UI:g(W)I]T,=Q
Ob]\;=Me_>Pa3_]TC,4H-AW4/R1aVe7LQU[FKQ/22UR0,+Wb0LFE,3+,G;3@S8EF
(fW;>6Id[;fSH8&Ib\4W7CS4g960P[RXdaD[cP;&6Qe/I><RK&-X&+T/d.9_L_CT
<L//0]<X6/H,--&^OK1D1;TKAR,[-5e=f,#>M3Xf6YM=:7]-);V\N_>)Ib#gG+WV
-dGBe^S2a_QMZW\J)VL]+02@\>@X]SbL<GbEdHI>F#M]HJ)61ND#G(IDV_W(RH0C
F5cG&gLCe:,^^P)bY;4I+-/3(_]bJ]AM>(>=ef8DS]Ib@Zf#<4cKR5R?6G9ES3-F
cT9_2&;&<<QK\BKRfK]-EK=1,4b_0G89,@S8WHg6^4MU8M1?:>^T/,19>CCZJ-D?
.\OcX?W;+DO545-g+(45SeRgPD0[BeWb_1FDY3OUU3H.D&^CDQ4JPBS2M,;Y^e.C
+D9CG]<gVb#L,.Y8aB3>[8@Y]EPO_F^7@FK6_M/437HKRdY?P#SD#NV8Z=@3Ke;H
#BV>4<eF4#+JM_YJO::#9b6a]^EAOYI97DNZ0aP7S)KB9QOKQ]7OE#^Jce<7;)0,
-Qe6c37YH2;K_KF5cRH+7Ka&JL#&S0U+L9=R>,=P\S.cL<eg9.DB8M6?Ra>9e5e\
BET(H]d:O9>_K5N<R+T,?IXK4g\:B#?C\I,-9H2[K&>0#.;)()BF0dXNDFV]8M39
dKK:2IHM>5WNZF8R-0P\UQ\L:5;bN.<^f:D_d-AUMc&bG&4]SbE@?X];7-)-<:44
Z#L>MDeI07XSbH-I8N#\DX#08?.6g&Z>NZL<PKV>/1Ja@4Q4E^)H[6X7;=-RZ7U=
g]=C^a@d&/06,H.ORKEg_ETWRGeC#=_aFT]f@TWSdaAM[,^5I3R[WF#0A-HFJb,\
D&fFgAW+#]#NSY8G86_,LecOHR<VaB7[NV&<=[UDfRW9.^;Qe\3(N+NE>0\BeH\0
)4UgG9/T2-PA@XRH2)d3\5H7QA.E=2C+V92WF6I9U_2MUFWJe)+6OPZ3)HHAe(?X
B;O6Z<X@DcFRRA^g_1;.Tfgdf#+^0]HYTU6:1]N2)-13X6&cXfC(6HVBL=3VJ(MX
aZ=E(YFaL7INNIF3;@;ACU_S_KQOcMBF,I8QfbJ4g-3Ae88QHIgF7.0a^+3G>+]S
Lf&Gd3YZCa5)Z/[/Bab=-V@ZgKNgAb0Y#QKag_Z0c/V;8-VJDSH)3HO;V]3)OS1@
:+^C9b/T>SICTbN=,e43G##K+g:F2[,8_Z.7BH&LN7KGLIH^WV7gJ7-YUYX61#D/
._;cW]+bY7-#ee<8._J^<b>.._;f4N2T[T3a;:A7Zg9e8f=RW=JSWYUGUE?c./\8
^]C[XLGB0W],Vb/F6X.g(#LO@I-2_2)=\fVF[\YEad<dA.])^)3bH12;+BYZ&(3N
0Q/ZJf;RLBdKX#8/-5caZ=>I?b/PE+X/]SE<6Yd6#,gP(5:RVQ-TDME;b]bL9Z(O
&3#<7[K+c_d5H&VF)>>/]#5(LN[R3<LMZ\2U&bK]+TQ:QAQbTNS7f57>(TII-8?S
G4+0.=Z3g36CMUQ3IDdbV^PN-@G34FPS9B1fA(&G3]&d@S?B=S>Y@K[Z(<V^DKI_
gE4PR0PJ,I8d_Y<8\+5f?=;&F+]D)I<<]X4cbED^K-\@Y)8RZU.W^b0FaZ2Q-&eb
&IJ:b#JES4/fZU[C:<B]_VI7(2g\FdF_7]5K->DSH)I(N#dA/Xd=YE0g.GJS+--0
961R=U;II#_XRTcUOB;a])EfJd&fJ]^f7JSc5<=L:a8;GFJV7Ob&,Q[++Y^0@54b
II;]^[21I(.UYO#:M2bZ/7A=STB6T<;BR3#(?bf[+d2J,4;LU0K<0HQ)XR.2dUdV
@bL3RcVCeBEK6#@@O+KcZ\bgTH>925_IOc7D6N8HP.G)VfUS7ZOYbgP5\8XES81C
a4LG-.8F^&.QF];01;8KZXCV4Y@].1L)RTD54L_-;5@?RGZa9d>]gf(ILHaXF@>B
I#JG]3DK&2HT(=]8O3@f>@IgD0^+ad+3404@Q]?LM)Af3B.TG:(UUaN.cK1#)gUH
JVY(8\T=CG+YZZTCE#]Q/aT-GcH/5QPIZ=@,,1e:;?B-TdCEN>V:L3H[T]5J=L0P
_1-+.3A9./7OHU[e@HEd8AB>Hf-6V&EBUFE&AVG?e_1.J[#6.?f3C.[.LI_CK(de
]K39cYX#=a/W,-A(dad0-B=^e#ASDA3XC7Ef.&WZdXB&L+S<fN9@#76@bP_[XfXB
g>:Ma>4ED+>)b[H?TfBA//V^R)a-7/>^U@]Ug-(UW&@S995)?)=9WM24Nf,?gZKH
N\F\<dX0@V2&K:Q[G/2:JI/g>,e;L07V/2QbACggF,0L;PTUO3OM,PA0d975C^_g
_6U1a3:DGJPdb_#^I6I](?X0eC2B7>65YT:<)R5@RW??_LZ,Y,FSe=JGOY(F<g@1
R=XF=&&2J<I,L.F-d6)0LO8-_5c:X&UcDSL+XJbK\U?3YN1?dIDI:&eB,[\OLIea
&LUOgY<_d/(.&UVZZO._0@3)>T85MWafY@;IbA)>f4MT]8E,3@HZOMHU?6gL<U9H
H.1H(fL##(/2V?-W7^f;QB0WO9B)_dSP?5L11;HU\<:=gRZbPC(_Q_TefgJN=@XP
@-==UKf^I96Xg4IJ&CBEL&g5be19JJ/b[E]3bf9[_L@W4eLE1:6C=[/<;YfQdSC-
X]K==FgYZgBM,cQV[1T5bbTa8Q^-J7<e[3CA6HZbK3cU&6?+^\<EaAB(97,,BE,4
A1Uf.:PSYO5^IRLHE^UNf<ZgUK[V9A-K\:=D;6RYAc9S_>6MFD3)e3HQ4+e0WURD
TD78LK;SYTD_F+:+[)4@I54H&V4eDOEX8KB_D.3)),]Pc6#?NFg1ZDNY8I@=f[H&
Z.SVa?@@86NX;<e;,a-@\\5Z.RfO_F)eOIa.VUI>D=#6LS#EXS#JUaQ;)-V4&LQ4
N>MdTT@.BPaU6WIg@C<(6,e./fP-\eB\AJF=)/DZNU,#eIFU\=PXd:NcOE2#7[N3
>WQdb</DC]I5=&bNE:RgESEgVN:CTa,7K&Q5AeC62?/7;F(,CIWX5d7?+?QcQ-1a
I>PK9T2;C?:4OQC0+E,-/=5[:7<T&5#L&YWIC(,NKA::\5YSEf6HZ[Ve:WH3+d&-
0U<X::^Y#gA,G2)0SQBA]0:GLX7PYQ9&8BK<);6/38&)P3,bBG7LX[#29#+XTIGN
eH5Ig^ga/Q,Hfa#Y:(]3,WE5PGQ7):YCLG8+,IDFK9INH,YONLf&R\dD.WM<2O/5
P7;@aB&[]-U[,>_R73/V6GESC_GN#L+dJ4a7DMf)OgXSAHV]AJAVOGEMY\8TVOUD
M/.UX)cW&JE;f;#=-aD]/#Y#SA)^#&5>>ZJ@5-QZI,V.Z?S<eaOQd_;_b:-&R+Da
gMRS/=?#99UBF+LU5OC\3?7_0)Lf9.+dfY7:#/ZO@4?MT14\8URe[:?Z4NZG2SHX
a6>ETRa1B+F:e9-B8g;QHHL?5I(PO_O?/,-3Y(0D/PU\\5../LaC.>&cbQVV(KER
A_09c7&G).,Za,/-.UR[\R;_T/8./(CQ>O&0OL[F5TA1b(]MZBT^@+Q9eX;c6c0]
R+gT_5-(ZJcO<Eg_50?=9J\>L0)5/NC)RZK?9adfW8Y(EUT(cH8K3&V:T<YOP66R
-LDfZFGfWH#gX596VB_WGWZM7^]6T?0-@N^C5/6KC/<HYO#@aNHWdXAGK?fWPI75
8G3D;>6TBKR>+GR6B-/JV#CD/Z)Q\_@RbKO2Hc<AETH\&K5GUOCaZTX5)&Qf3^Ad
+KUO]U,c:,(^\5e(^P-V/CLODQ/.;,Zf8M&LYX3eaffF5L24T-V=J4g=6ge4aXV_
;8=+.XFH)<dSD8OWAXTXb^fC062)<5@DZ]+ZO\.JgA3.9;0J_1(CT:)P7g#N.20W
#[863<B+V&3HN35\UAb:#6F=<bSH9dU&=6LW#5K],eRV0#SfAS+9@A833=Hb(MbD
]DOFJQ)GQ#<c.5^MdPQXW+6IN4M:_4/YPVBXN+Y.C#3?3\RD)JDe^.=#EBY]G(9>
RI?bg5?gf)EJ0XRV^-@1c?g_:20_f/@?D_T-#gP,Q9AUWe+:OQd<L5#F3:S,DHW=
[H&EWXXKK?EH^I_T3=Rc?bRL82+FV&^7<\OeGefG8GHAgE=(IW9#4JaU/2FgQf\Z
>UI]<[H;RQfN=E9Ng33NWL93:X;.Q3DQf2CW6C8:8,+UO1Fa)POG82PH<fHDZ-YB
9/G4Q-#UCPWef])OYNgJPX=LY.<QP7JWD>CWYE6e_QN/\3:KOZ^&e<[)53N5I-,]
^1C,EO-1H>JP;,#1QP18(e3NHKA=de[@IfIdPP0Y@F07A<F>J[:c.>NLfecfQ@>B
.Q@017G)3bb434AYX+VW0IFAaM5<KN@d.I&U:P\01D:R@9#57cA7:5eTe4=)XR[/
a^,YQ]+bIC#D7[6[Q0:DTHa09H_aR^+EGcT[TOQ&^:OdFdW\g(T^?902)PdaJA1:
5<4SW.CYcS&/2;]N,WFUJdc,2=XW-;gL#KBQ-CK3KD^R#I(#3KD3017[Mg[=edd\
b<8g>A:H.OF9^@-aN:LaQPRfVf\NYNRO0U;5?\/P];R69FAN7/aaD&cK._+X)C^1
C:Af.,YOVX#Y-[@\LNgAI&gdX8b59(5PR:@B?-MX0B_<E(<MM[RLGGV,-@@@#D8N
/[We9M(Qa#NN<LT;4@I>O;F.#=7X_VDYK@U[M4YAST:VDU7.#/>Ved4?SE:5;d)I
]aST0gKM,3;0dR@0MMGZ?2K,>gM#LgTJW,f)2A:@=9]+fADG1\aE6K15YP4[-1K/
6,fS57)T@&C8=6^Qa92-/7?938H1YcVLLEY4-?<6FZ_,EU^0IV;E;e0U)(U;90=A
c@YIAQHPBW:.,9C7KP[JGJb5EaX5QgW+U0ESH\70(ZF?C)bKgSe_VF7>4UEV6^Hc
2BJcFbf@-XI<eX9,X6be;+1T=[B3]WHYbDNTFHZO3[=?VJVBJ.-?@W]f1)LR^S\7
?2NFH(?N[G9UFNd<+=X0T4fFY5fR?YHe?B_+SQ\J#?ZcV;JbRE0=V?4B+WP>QWW+
XPaT=9X8.XOKc1NdK,@8OfAR]VbU#Z9N4>1[_V5I6NDJFO<F:MMPUZXG<)QTA5A&
K?,5eRIecRE<(?VTZS\M8bg]F-0+LG]SC(]2[^88,DAa14bSFK;CbLcW-1V&29^-
abUA=BF/4RD<4HAI,e>A-1Md[(,?Lgd7#-7X4d0\EOO67DcJE43CddEE#TAD3-D-
/6&?JRQ=I4/5#@)W?eg47K.^9Z^XIg1M]P6d(+aX&K&&R]/IX[&/SX0<b<D3D>92
AEK2N77[QJA6Z7G?0&4d=&@5LR<b4V-3C+6[>V4IQad;\6TcfKONFY<N<g<K8[H)
(<\CV:Me6Q9I)B2DQ87X#\M4;L==[=3.fAI=?1UB:=0[?F/d_BI;&gb,bTT>GfOV
cbcIXTYSUHf+>1/e4S@OX?&+-[,8I?B,Z74Re:9&aU#?4L;e,])QGA828bP9QG<R
LG=c=2OZ&1<S&\+SK:1\+a?(SOKS&Pg1;,11/.P#MFSg)@NDOG@<Id(:PF-P9=#e
BcAd6S(6M21UL?.X.@&dXOK<05W#DX.)cJMCHEb8FL::/O8a_V&J9f1TA^5aXM^R
aB,(K@IeIY,7;[UY^3)Qg2,Baf=YT-9I1M>N4.O=a<PJ0]U4&EXg<\YDF:LGSPPF
XJTGVU8>,]GYe1R]8K.6S8?,d#Qd3NE/&HgHgYgI]f<KcVO_^IY6a(Y/22-?:Eg/
>==+14(aI>>P9UZ&]4JW[Q][LLK(38L:S93b\K73\Q0W5[U?_b3NUZS2FRD)Z^dA
2HAF5EISG#:P/:R5,N_OEWV.V#O?:WdUA^;G2UAQP0O\-06UPN/O,IP<^<]dK,Jg
^f0MGESY1CUM=GW.YR8]BJ?;>,^AV59T9(N<3)N_<8^]#?S^2V.R;/&GXA-O:WGU
U.K-JTIcWIG;L0+Q2RZd@N2)\ERYVQ\f4IJO-KCHL\G<0JUP<V<NdQ:NBEE/<Z#V
UaU]9e03+a/822d28Qd)d4-R<Z5:TE-&[ZO51\@?-5.5.&,g?D>D86O.TPMP.9RC
VD)X&5DMbU6aTD#TP@\]M?BYRaa5:gUSdeJXYebO9B^Za1a),8#4\0)P/]KKYI7b
d0@B8>Y)G_+N3RD,<eO8)=@T;LNQBSG]ONS5g00&W&\d>.PI2b-P.WM&Jc5+P<J;
<F;4V-,6B_GFIL^V/I=Hf&TF/G\[\NJMbWT[N:/E:9\e4I3J:X_^L&K#4:PA,<^N
ED@^bAQ\5]X(;?9M^+c?3^(D#<S1=ETG8,^VW)E7N/I#TPL2Z.=PSIbYR&[D4G7W
KOG2@0N,,P0bbR=R+Kc8;NI)U#I-.G+US9g\NLfH4]e[#GTaDD\7YZTRe(\MMg<c
eI]@,[<:VEV=_EG&bB_@B9b>?0Da#D7(8b74gY8TX(.b;3GI.G39IO-\>PReb=9@
XEQQY)\;5F39&Q.8[?XV0Hf8UGO1\(Ic3P0a1RZB5CPD/V+=V849TQBAQ<J,:]C9
bEHZSMP>FXA4OT14c4@KG;N)=bAEGT+#JH9fce5\D8Y/^C?Baa>]2b64/g6bBBJ6
A4;d3a0[X#TP=;=;]AS7Tf60.Q_^/OI0&,[f1Nb[MPc;QRfC-)SR_B_\.2SPL.5g
<6VHe&@cSO:+L\_B07FI+LV1e3QU7JN6A)A7:];01XG_]8^>QM.>]0aOdCF\Y0QJ
N[K&I(7R2_Tc]J@139QWU6GF]=CRA8_6RdgcXGQMa_,EY<M<g,BIZ82&,#R@H8Pb
c-:Kb8HLUDaV[>a\>&^^=F)/NFEWG);LVD4DCBFJU</Ya\=IE6K@b[b>DOdW&@>Q
_DPEQ=eY(PD#B0.:Ea^L6:3\K1[?2:U<P4ReW7]#38FSe_f+S7&2b^Z2@:QE7.38
&WX>6QIO=H.(W2JXMF?M@_1AKB62[]F-5>^UC_M]N@9?8Jg-&E;39R<cKV(CXPZg
)VG8K,K1NJXON\<R49,@Ce2g[POA[O<c?[bIGRfBLDf;<Yc<P,G5EAdX;L4MA0[:
_f./I--gH#;^bN&\bfE24)6O;gY4]V8@?Q:W-;2,)#A5eM,gQ_Lc#/+(^=6@R7D.
eVNSCIVIgU)g/F9[4.DLY;0I)QS^4B53c[#,2#Je_4^Ac5XM>@cAE^<8+0Oebg?b
5PZ.TR5\Ee4)QL)X\,9Te4b?aDe7<BXT1f>QgKM\\<=0J8G/<9ZV.H;]+6+72VI:
:/XeILRW2B@c09ZS]4++@>QU4FB-1S-;d+K@<&84VN@K&V/F;@S@8#<G@==16P73
:c]K>;]^eX;g8T;OgQ9-g23+fO>-3J11IR\&H5#>ZU#.7MQ7D6g[5Z#3=VX8dJQc
I./>,LYd9Z^)U9O\g6>eaT+,O]eJ9B\7<O8Xa9K3&#,Mcg)8c3.BB._Y](8;HLNM
e3^UU4G-H4O1.#M\<[/?f=VHKNcC>K&9^bZOceeL5]-E.SKAYUR&C1Dg3Y>bLQ_<
UVRIO:bC/#6e)]b.\_Y5d>d^:[=-7<TC^HD..CgR3TfTTPS_g^[)7^BV;\K)e\Y_
CK?0[-&11Q,f0EZ1eOaeQDKc8[C+N]4-IJ)cR_..9.#=YS2Xg27Ne&XONbGCP-;c
Bed;7WN5bINKTBa/:337dWE:UO<g1)YA:CdGBU4[^],SfZ.0D.C?V<7gPGTG/I)<
RH@09]Qg^7DSeO4+7A(dP?0?]_@:8ce/C\ADQ]7fZ1Mc0+-f-H_G6\)25bS)BSS4
,\.:6FX=-S;0.Gg=M]#eT9;P]PHDG0,G;7&QJ1,W_5)ObE2SZYIZM?+^3YHC6#D<
R4d+@+BeFa7e#:8^P82CU[@MK/[^3I\Jd^(f\K10A9TJbP,Gc(WTS6dEV7B=(cY[
9=]M\^c7D<D,R:N0F7V-O=dK.L2_EBg#PH7M73fC=_d-<eBY_-?=@KR&,<@5S\MI
fI8.bCe]P4&2aO&#:C6/E<CU^-O0GB0HS[UWMZ8.^D=.78K,AV_@.E^7e9]]R3,/
A=g67_;HW6d9Wf(L;J5Q<<T5G-Q_g#/AQ]Ze:\/DW\cKJU9MLS-;;43+0g(d,I98
)Z=33C^8NJHE2fI(WW4^2NK&LQZ.SL9IS1+3<0Ca#0DbG2HbSF]<dA=6Bf<^)PP]
<;F;,#/R-)gN[GU]L<_6c4[Q;HdQO=ZT5(E6T2dGeY..Y-_6=GgCA-_D]S6#0M)J
EQa9TC)VZ\fZI6eBcGF,39KP[P2TS,,Y?3[6#2F<>)Y[_Va^4,]2.5O(DD[6CY+H
(95Y&<CaZ#e4aJF8(9C<]AAZSVd]9<?,\6BB3I[?2eX9RCQRVcHU>.cD,A0^^<\d
6.^Ha8bT1GRaNGcMc4bU9[5Ua;???K#aC_&gLQXd51(B64T)(<[6S9#@SZgEecG=
DS_Q-RAOIDOFZfBN@F1\TU+@Cd[@TL=/)cPS)V,a]dHT+eC+C.gZ0g&W#NN770<3
g\=2CE)g=JV9X.1f@Sc3ZU@f#ZW\>BF\JX<\@Oe1M[BQYC=.AEZ-R._1=#e\>aK<
;Q1([DgE__dB5[Xd/M\)b/D?;[DJ5.AX0_P<dV+X^2bFf&4.MMf\H8?EMI-&CLLL
dLF\30TCVM)S\PK&O>g;I<;EC6]1UK.Y:<;=Q.<0\UU;2@ZRI:dW9>dS5P?eKHF:
P)?cP4F>g/cZTZNc8]#3_UAaE\,7P90WS>>DXKL-#PO,\FUVS0L\A4a>Z^QI.GI8
@NM.a)B3FDK++A<8[^YC&>9\@TZ6)@QUcdL4#\8\KAEC[S-,=N1DJfP-O([4>TDT
5L\.ES^VVf^KM[BBYZZdT6=H#4#.JIZ5P3X,62b)#ed+_Y\\O+W(Z0UfIM(Y6,c:
#3a53950SgfeM?5XX3PgL[d4ZD.)ZXVCdNSD(-Tf(&Y5cB\#_&</[^NLN)0@UAU.
c>=RE2aFfPF(?]K)5=&Je#\SG98eV8Q1G[]YO&0X2\[^)7FMU()K@25/SS:JV#c#
e[J<ODPT\_M4geIT88?g23CgUV&P3>9IYI]I_3>d9f0aZZSI@)DQNJA7=]g=7M9@
eM]I)V_b-+&NN&JX6]\cOQ@_a@7N,HZUgBcH<[N\+^fEbLEJT6\Wgg+:^&++2H_2
Z2E,#MVEF<CDQ0cAAF??PfT<b,+d0[=OUg]H=MDFD,7Y@gU,JUaa5]GK.B:@OB2E
NA78@Y4Q5C@/9]4FgC;7J08A5Q69cU+@M#=UDDVC<9<>T/eP9-A^1gUM]e5DJfJJ
c74Gd#P975ge)<0LG:2JW:a<;?g8JM;T(C=/=Gc>G00+U=O7#g8)C^6-HT_KQH7I
b2H;F)4eC63YSF9B.=.(YCLE9eOY;927MTO05#]^:,FS)?B5GNH6K237TF9#Y9^8
X,WH--?abUbBTKBEf,<F40W[b8C&7)S285C>3V?ICD_V>_GP:EXLB#T<fQNJgg?2
#C6LbD,U:(H&)BYT3g<XI?g/USKd;2O/>b=LK.F@Lg1FK.>_LJOB:9Oca]M\K^5f
[WGa[6)-H6@M,CXf4U(2b&UVM_0(3-D7VW@=X7VVce[C,NF<Sg&&M&0a/81GD&d8
X/ACE[&[\8YPM66d(B/63WIE?ICJc#MAK)2)b+^?764KL(D)([:ZGd\E,E=#=H[>
1\M2O17EcZ^Kb(f=,/2240@RG,5BBC1Kf\_&07+C6E;[2b&U#E99\5gXM:^^IR,F
K:,:IJV5W)TA-ODQ+6?BI;Eb3I19ZTTM74+0ac(:KC<1LdJ=5MP?HM7YG[#I:&X(
)<Rb,X?:K[>9fEdW_K]JJDeT5NBc<?OX[@bX6;X08FCJD.-C^:=Q;]QeT2V;YKVP
UL2XHc@fKWP5/aAQ5/@C0GfSQ@[56c#V<M3Y7b]M9EgW@Z5TK6Gb.M2(&X][_beT
56DZ/)c9E4+64^c>IMSZZ8Xda?[X9I[?>+.U.O_?XT-=SIBQ0OZXYEJGKcXR=d(.
WKYgg6TPYd2=>);.\GH/)e3:>:+F[82,+C3W92g<2gB(5#^\IUeIQOd[61YAU_f:
/JGd=D4F^dB<4RM:E-F[HW481,L&JT[1\@#Ya.^,d27]&ea6^70M/4)TBR>X>29b
K(&:\NL_1cdEQV>^6;:CME]Y7\0Tbc&90H,Q]G2A2D5X7L067#QVHJf>B@(+M:ME
-f;FKZAgA&gG]GD-7[7EB.L5G^=/+HXaNY>TV^L4R(ZPSc+Q:818>-JQ0TK1<3+5
I]\-2-@-fP]a=>OO>@aFH)U\1b2;@S]Q+O6g]/DcP0TH:,aa;C55#IV@RY=5RDJX
V9LGZb0f,LWT\(fRS[41A&>_)K8AN@0S4LcS0TNZcM.EO<#.-H>70#G3(+>eB?Nd
RGWLZ]c:#AU=O/UfY9Mg/45PL;c<7^Q=9dJ]B-);PUM0F(+NH/D>dZD61;C.PH]N
-;T.?QcK3;5(=A2]#U/XeLDd>=,Z<M4)e?V>NfdQ4Q]?D0;#)F1-C49?40^Y,Wc.
8@0)?W1<GDY;-<A#e-d(_JT,3P5T=DNC5CQFc/5IO9d45-._Tec7A;FYLFd1A[d?
(e^3D0bM-KJ+\:&LY;VdaN:R1Z_E\XICPG6:#.JGWVOVK)JN#-6MJ0gGVN08Lc#:
I(Tb26Eb.^a3:-Xde+ETEf8M@9M842QDMC/B8PTJ(&;U+A#H7f@=e47Kg5ebNKMM
0M[8F<T550F4aS?R58Y_+,GS.D5#&TO\G/d.&W[SAR&5N#J>)4G]E.,?J7.V//5?
BWc/WaScRFT0>YX4R:TX&3#<V&_f]^A@7LOe:OC::Hg=AbfQ+_[Z;-DXXf#L:=;:
aZa5W,SM8N6-46_RLF5/Y+HP[CW65DM5.,1RHDVFg;bT3Gf8WBGF(V#;?-R.L[@)
U.beF23:ReG4>(d2TN4G0dU]J2JD0_\aN8Xd1eS(g])b,^WAO@H;J:<53&cB]14U
?8O<&AM;/<C=?DBZfQNGf3>Q6KT3FcLMeQP,YOg:?D^[6;@8RCAY)D4F6,BMVd7+
=(<TK#)>7PcC[+@8L:e57;F6=4b2IQQ8c31e:dc?O0+74K4+W/Yd)@0:6W_>P/,Q
6Qg)YG;X.;U/._@?R92dg#S;:OZQCfQE8WFVI<,]RcWD9&WN8MDIe\:6fO=T/XR:
@XDN1T0;&QG^8M#(dK^a(Ye;?d?)KR_Y73]^,Q#0#>)e?@c/SS5=FUV,ZR&8HXOM
2)LW^N2/,_C3cQU9@:Oa_A6DLCeI9M/Yf#gaL&,D__b5J><V0V]+N9)(QaEg+e/)
J8.S@#Fbfdf?_,1>2+3GZ.@C>.&M-_Z3N>g;B(J__Z]3_-/ER)PdZFW@VTfS4/H<
7YL,Q?(58A]bP-PM(+NWd_c238a##CcWR^/9Cb)U7NX;_N?b6GCN<c0d;A.c[BY^
36B#O<]O9-+L?WG8ee?OCY_J/_>NX,:,+8CUZ1&Q9bPP,dZdVcWcAe1#CMZ^C.1K
dPZ[bVL95OC;:<:dS@]GXA-]>_W632aEAc)[;(]N/7DI1g00^WY3Feg/Q/=K2GbX
\AFQ9TG?eT7P=c]fMW<EYUU\D)e8Od8eH[7OQeSc@(UZU.#gFbJf2OP&OQYaCZcN
&ef2MC0Qe-9?U@=PD06^g[,CgO].Y9fb]A(R\43TH(WMO5<6+MJaD+-:270M#URB
;8@TZB21W^ZM=SIL[FNE]F[DAgRa7[\5AF2YVLW,:BVBZL>]6Fa&8G[A[A<1Dbe<
bY2;:7abRK[HY]4#g6;Y:G+d[eIW>U^_dJb;C7I#/U-LcYIdE@fC#Ya>VB_##(FC
HHGSB[.eX:NeW8=ER<.WHFDC;d=/:ZHC=6=DBJ9VX5IVI&P[482+Q7:7P4:=R3WS
:3YYMH\.c1&98+/b=@@gEAHR-G1:T0I9A(Ha:BH?RA\,)6H>?/P/K)WVJ7a;cO;#
N+_eH]HGMOG@#XDF0[83V3<(((Q&1OE[P/+:<_TFH6Fg)PN2/J+ZO?#,CHR@R]?a
3IadF:Ag<Q,F>EdM)]c);HJKd5211RO99]3Pf<_^NcD-/AQYN5B5eTHe^#P/?dWS
]0B@ADC0c=:aR4(G/.[EB,W/\bKLH_+e3/LB:6ff)83eTC.6O9_1A,e7U:DbUP)=
QQO61gE9)?NJG06GTYST9V.CI-W.X8T[X>aW>2MH46]Ed1SEEc4]NSDJ0Z_NDB9C
cS#CRTgZZ9cFc60.X^da-GE>eBAJb/Af9ZeKREB#:K42YMbL^5NO,?,Y-Q7:(;S_
5>O9-8;5DCES=]:ETJOF_EW,,K&;;a#P?9B_]B+F1(BTHDd@#dCXRdSL<LMdSQ,a
,2A<G=GN4bN;,a5>@K;N&:)^f42fL9-<\Fd[D>EW@;51(aWbRXOJ1b=(8+VE2e)<
X)&]Ld1+ER.?8.a1_YdQ,_G5ZA0bg23A);:1f?U0L9c.1a2<e@2T^;&CNXPD9G:5
859Ud[BDYZCQ#S.(V.#-\-6_/2F?-NBB>34FGNT_E19_,A_1F,)Od2<U7a_UgN=D
3Z8FHS4RMEOUeAH?.08FSF>a1RJ2_Q-+9ZZA_&-8;ZZ7+31CUO;W;N,,801,MB4C
LYT=:X[&MJHB@^4_bAb6.a06\YGW3@#]dN5fJ/.S\6X)WGK=<(\)gN_-#+MNS?RW
2Z,a:\IQ.eP^^9)MP><H2d>bLV\7:^C,OcJNN)5\<f/1=@8Oc,_UTL:/d,_&DC]E
7)_f,)GXU+ZB?49Z3088WaITH/((;(d;]090GJ6D\F,^PWRL.)E=H.[VdX9d9HAe
+/38BcF#NJ:FHfQ<.5;HU]EFDIPGd<AE>1AK-bXDfM:I9Ne.RP^\HSCU>3_&BP@C
b#&.#gI;,_ZSW6YGU\SABN6KMg/L_B.a4+)bA_[bTA@)-56#OE#<S>51bJYJ]>(M
;cUc3fU74#Ga)YT7b+T)&f.OUI+JGT+TaDQ)=4cP283eKE.9TEK?O.6-W,AIcK&W
&8D,GabMSUVe.aa3gP[-62B0.a_)K68:eHa?\OcZF[V-D5]OfZ,-[B4[VA0B@CV@
gVK0R@1VeU_L6)CI4)8?QB#\;fG,)N3CHRA7@THZVe/G^?;8+G/dP88H;L65_-f<
EG-@>+:eJX:1=8QX1[UC[WTXLOF34R&\1ATWASR@]YWRIOE@AOP:([D-2IV.CD1X
:4Y..V,]e2IfC?PI^/b7\>GZ:DIK+EH]XYJ@OJLG<+e-d95>Z@FBZVaUc0190TaE
XWY&0XALKLJ-UCW[+bOD?J.79c61/>?W=.[59Gg926Yf(AJ?M2CG?)M&0-.;=6C?
7ObK,&2a&-(&6dc6\6KE_A_^XPfM2VgY0#d1KT[=HIV8X#6L7eDg//Q<^>]..Wg-
>Y:V/)^6.?7/K9SWY4#EBK8H29FJP]3/aZW5T]\:-2:OH4HL#2CPC5b_NM-aC388
H/6)ggU,cd)aY[IZVOTY^4+1ED@[]WUHacTeR7Q<R.Q-DbgWY7;dJ9:b/cdJIaK:
.2RF8RQ9YPbaO3?X1T@3MNZ,eEaQ]Pf2>=88QK.[:LER?#/_g/ef<Y-Q3)R9LJ;C
9G#D3g3R,g^S-AX=#-3^P97NEgbd9,@^]D<XM3bg4+J17+1e[I0G=9cc7RI9Y^c(
7?Z<QXHR.a?GE^\:K4?P\IaV:OFP@3Y5Id0(D>cQ4cfS2>&+<#79H2PS[0RWJdfH
f-Z[L5_f&QVS&g5Ra\V6ELVD\@:F0BdYK]?8U6C>LQc9CNNTJSHX\.@Wc#W(?DSM
:-\D-++5EN,0\=WcGDO6d35?,O774eb2[)Ca.^]F-VY5WPP:Mf5;RX(,_(0Ea>VF
>7N(A-B)]e:,O-1;b]6Y?#5+(^-?JF9OQ)J/M=gS/K=&0;\F\#MC^J4Pb@UPLUaX
bYX3#NG-Z89;#CV7,1?>cNWNML2>S;UZ4U:+?_+;K0.G-1bL_C;#FTA:fI(I/OPg
XZ\:YcB.1c6NaNgB_J#BX7HM2T2#_-g:24[.aU:3U>DC5006RMUU4KIRWIb[NXV.
U@:EcTKYNFe7RV//(\1#I2;_gg;Jf,V/\<N#G&J4I@A;c8FN00c[,WN&0e7M?PK#
SJW<F1bL7\1=W#-O^0a_X7C_E4e2T]d?:LWfF7[+Xg0^;Kd:CW:5f0d-0);IGSMW
U<5-GL[741]2LQaeJSUZWB>Hd\8AY0+JH)-^fCT/8fZSCJP-)ON#g\&T_a;a:RF>
9:<2-EN0.6I8U/]D]I\]NbD1I,?;T2^:AZ]X;\CLCcXF[GY(D]CWd<N0ER#c9^0O
=edYGdQRd3H/M].(/(<<G^XN[+8WE0K2\BOI9D\SJ?DYU4KUg..E.V<B>_#/F:NB
B&@gJ:dB.XUf3Df;9.HLB/\\KK.MaZa+d4a\KaEWAaR9Z3:f@=FfR)?;&RPAN#4b
DT]CFA0QW#.G2GX8ZQS:WJ-^=\e9b-5=R0D96A.eF96BP.c.DNd(dK#:/@-R6/49
@U2Yg=/6dd/,8<I;?I.S(D9SQ:HV.A.Ge0Uc^E>_PUB([Sc9e^_M]-JC=9EK?GM5
_WH,]3SMLSb/RO&c)EMfABYK&)R(=c,9e/c04M/+LO\FMK?--J11.:0_0VR(M[:c
EQ2/(&+aJDOCU&4+V5.O)Y(/g#(4.ZAcG9_,6>QH8FJSWJF1T?M([SK</#Xf18Fg
NeP;\1a_@O&0.B;:>9O<_cML4_Z;N(DXRIVH6ZLMAQ\_f]\Rda5DQ8R_?=bCZG_f
RSS;d<W>@X=3S7=+V55E/J\Xd3D=@ddf)==;O\U61dN0BVTf[7A@SQ?STA^P.6;L
9UHV8bD4&>_.[.NAPD+[R,8QPRE<g5WQgH)f5IR?@-AABECIFZ0:;-[V^R:8-b]V
I+JB\F8W@#UQ@PF^Ke[OQS+6G&TXKYODb;HTI;Y=.4;FD1_9B7<+HV[AV5/LX?+6
7:ga?;1d1.2W+FGF<,B4G#LD&7[MaM,:\8&V&&TF,>/4YJZ0Z?61Hgd&[<eR5NZ)
9/cC?PO<+@0DSb^IcV7cXdA#.[TEC2<IVWO[SaY/cO^:d-5(aU,X>\N6<fJAA0I9
_bV(eH[[EKa_D+AZ0A@K^SX#&+&HS,c#XMY0+L42gL5IGW_CE==fB9ND/d;d>bRX
/EBTA23abRf0\5Xc3/MJWO_ZZgNeO]1N@9:FTZICS.77eZ@&V:@RW?>RYEI3W)ZW
>f_c>M<-eDRa.[),C9QBI<Wc9A0:T3)LH@_e5+D=LCPW^+Ba?\8TAJSe,U#HD=\B
BB:FD9E,R=3G?RMK2]8HcCP+IWM=eL2GPM@gc6&+Gc39cY02dJdF=aE1eGdE+Z#R
(;AU:>U&AeCXBJN_&IF)WcCFCX0PZGHBZbM4C.1+ZI86FG,bLA=?Wa6cF];CV7]V
>X,MH7b93:#MBLEVEggfUF4HZ9a\2^5Jb-WPRTdM0JUYNDbJ]^c(+&Y;;)bc@Q?Q
S07d<A:3d8R2aJ/4H7g:Fa6JZS@ZYT#@5MeMPKS?G<G7X3G3K0LWULU9_0?7[VcG
XITE&PT.Y4[YFMKH=@WP]UfVdV54cLH8^=)6KJ<?>0#:1>&K@SS;ESQ+ef2Jg.90
E)Z=KG,X1-IMWWBCa:bI7<=F#acB,BgZ92KZ34BPF0@VAA/BO0g)YcAUK1=cZ_M,
R6E_g_9,?3EI7>DbYKSA;\2e=YEfWV8:W.V^CETOUc\Z(_G9&;e/&</4H[S.RL-H
gGE^R#WFRE4.&(d.GE83NH18BUDMMKG\RN:0bT5F6dQQWN]1(4,+c1DCV\Pd:&D<
b[e]\L(4K<5YU9EQ9KH#MY&D;-;EGZ&\KI(VZB7ca_<+H1@<(;G#]RB:;?NM8;L]
B+>L&^J^d?-GOKS6[.4O=YTR(#Y/2MI&XWQM8)M,>fVTbU2D+<e-VM6ZD@.2>Db,
[B.:HQLAY-b;(KEGH_S5RNJKTMb46US96VB54TU/0FH5-5bLKIe&5)\)>IGG.8.H
>/I0@d,TCTf#U=-gFf,Z_Ic9+6QFS/:C#ONO5=J,X(^:[MOW73O.;1S:A)<([M)J
S+[3ST0F-YZP5&]1L+\8g39#Sc0GTd;Ne]W@O-BILA9N/AI)/a:1FIK;E9;7DK0E
Ag=RYHaU@#(QHME+BY<TYgKE)4_Rf4/a#E&&8NECQFFV&-P.O;#X.?>_H@-gbG?b
EYMa35Je=dJ2c^dU#R@8\We,Hc2?HS(0[M5#TAgA(@3))9dS@gI:cQ#JOd)E(^3S
0OPE[QOKb<f42J7_\WIHC\c]J?acCQ/(b7EEPUA^2&KIRc>>3MOWJ\;f&^ZKH<JV
^L/7eS-MW&>>9/^>#F23,?eXa9N9eHf=>^_3@W;GYZ?[?:eBPcTb=c6b0)>EbSW:
/:_7#Ud8(g[OR_4OJ,PD\VRZ?YRT7>X0,[/f1G(GY61N\1CQd7+KKgV=L&T-9/62
_-5N#W/V^C#\&XS/+5HJ5a<J(fU8WW-K@)YBH.e+3=L_&>:5.Y(e_@,YP-042>Ya
[;=Y;b>V&GOL](>(U9[K\(]F4cC]=ZY0d3Ia8e:51;<RE-S_2[<#GWK9Sg]EO?5E
LPJLcFN^<)61.ZJ=aGTYfP(CUaRFf^J?>26>gJDUJ&NF9V>+JBDT;R.:&KI\7IG;
3LdP(bfRPADF=dZI,/d:].>b1CU&0]+6\1RSN+NW<WK&YOBTW=Qd.S>UI^.IFCbb
.?HP)2&5<(I-GAdEJ>WWKLV\,D))>fE8-#CG/)R<_CdU8C=TgS?Q;?#.B;;:=I7K
T2>,)PGCY:G^UdZ^>.@/Y.SZ39Y.4SH#[(,R8B]NO-KXXc0=TL71_cJ@\eK=7NFd
IgS4[D].a>,J(+M=NCL1THHY[V0B9g1Ff.R9E<86D>)L@ALX+.D]bR(DTO.=;HSO
GP8KgZV0S=WXa9N(?W]I^6=RL(EVS2AN>-9OWVRaWaN3F1#0UQSE-LA[Z/^L9eOa
AI9B]MM68=RS@MgD_1(NNO-2YG-)^AA-SLTK;bO5-6^N+S6)+L:LI@_IJgU_OUX[
g_:K7BKBDK_GR,+GMNE)8I0df+b8AE)[,6M9T(].H:3-^R>aPH?#P)bc/HQ@-[^H
T]0,0McG0fgF8-]EUYS2>UMP5#-.-/9GQ+eZ0>QdY+b5XeE6c\I8==?a>7>F61ZE
AC:8c2aSPO5E=FAg=>+<Oa_G-=WM[&e[/K20&Wg[bg0;DYZ+U(DY2.bcUMPI<V;\
[#fWD(S_bIIDDQ&;)]_BeJHMD8f.I-R5^<EEC1#)XXFdDC_O?W(03@-dH+VU4^#K
7CRLg/7-_g>/CLP(L&,GSB#-1#)DA>TXbe,gX5(4C^@DfXKYb6?Qa=1&R[/L-9QV
V#eZ4=0ECFBA[ee1(&42SO2aX>C233(T^?^9&=0K_)B3,PeTe6<HAQ&N3E_U,f/&
R2.GYH9N6SIg,V0</),X96&f/V)EX9S.?1#H:P)7e#@g^8(5BRAdKBWDLa=e31eE
+:WMFCMBE_H#edCZceQ\0EL0e#HRYC\E2]UdN&U2GW(WD:#FT[E<\=UXT+V9f&G4
RB[5Z5K)3GVA=C([5>B,[:,W8)+Pdf4-QCJ)4R\e,U>IVC^.OP4CGa[GLUK],Q=A
,9+K:c)\A5A?gVPN[MB>&+8A\[8aU)CDNeVPQc0ZFg(/df^VH0b2H.TV8EZ#7,@0
U66UNcOQd4_a#7,PO3\:c8Ag9E,6[3[S\0OG=PAV0TC2=^D:M<]R(cc6a(TCg;@0
MQ(4HQRRKBF+J+VUK;DZB4X(+>>3^S\ebC24IXA=0O4WMK9\I/YGFV59@K:bg[gL
-YKK0LedY=UHB1H).QD&]LR@3()NE(F115VC(R3b1cff:->Q[cfAdH65/7WA>ECM
XRTZAegQL8X@a0KdCTB(g5DTMg-VDU;S>IJCB-^=0F1b@X98T>D=<EPBag7^T/-H
fLa1(gI-c16:d=4&ZCYI_(e1YE.ZCOB6BJe\E0-6@=1,S\Q4=NaLQ^BL.-8:cbYC
T\[H64GJDENa(3JId2#L0QAZ(VL(?<;3U/MBOZ[80D#e]<Df)JSFSMQ[O4Z7_U6=
W3?E9:#>;:7E\\9=?U57Zb-C1c;4T1U/)&D;>ce1/JWa2^<(STR?f3+LD:8N=/4\
Z5YV@==EUbJJE+P(W8HQe3ALK?Y3S<B_Y:FE6/CZQ?Cg-_[SFJG(E1YDM)6Kc>GD
L8=8A6=X\d7&U:C-YDI+G4#L).<Y13:6S7BH3ORJL;UC0EdfRbaga2-/g12b?7A<
8c+;]e:K0N&N<e=/ZR\da49J)1[S(+<eTV2c4Ke#TN1^2R]4WFJQ,Hc0CUSG2ZA1
#<gNQXf>A2T<=L_F>Z97]DU_9ZY^#76A(CBG-d\E]-&ZHL#Ye8];@bQRCX5]aVDL
8:9J&7&:H;MWQ#[.#S&>F-VA<6@LJR8GF9PN2_7<1[TR7gX?D7458Y4+IFYI0,aG
H<^(dU4V5STg(PE_>4K9AV(L42N3H#DXQE2H4BE;S@UD11FB@9RT9Q0<(^FQM[[0
TL&cH.^;Y7(c-@JWGZP)eV:=2#E#PHF3Feg6?0#=O4.3f8O939QBHMN,Qc:>/-(V
2Ud)GTBcR=>0\#9]P;DGJXB5BV/5H+([:Z\&-6JN7&#4][X0(7Id4=g62b/J_0FW
G0=b,YS1(]./[PAL[a9Rd0XbS5<W++;LQKbP0C8fPL\K#C#55LM9/7SX&ba,MNTC
EZR03#]3f)-T9fg=BHg3L9)]20:QHKX.2+PM.PT1SHM/PXQ&26/#6dTO,\,:/;N)
)4CTKdf8U#fLP?]5T9]e:@UJH[8XIVIc7H+_6@C&;E,F^1]PMQM.]fIUJ>f-E+Ya
5_>I65d/,,FQ&JMaEB-?L8PbQ3?DMU@JY&SOAZ0V7Y.)=Ga))FP2[W+L^:U]5-&1
[cQ:_Ufe]Z]?E&+Se/W]A12OBcaE1-(IgX2,_3>7^H8V7F5,7AM_LU0g^NX.L3[.
(0^-(+.7[<58,]I0F0R=ILWd.2R;7O[?\.fZU3WX(WO6YcfeQ[O1eOe/b><V,JTe
DWL/VR&:#)X7&EXL4W[\g/^[dM7CXT6SGb],=>\@Z/#,c-/Y1g^:OL8=Q]OfD5)O
8=Q8QJB)[;M\ZD0Q-B0MgHJ>;>5DM66&f8YgHD.cg-+2(IAc>V/#dcQWZ99HCSK;
E9\V#gY8+(L/T#<c0Z8-d>>/.5LEC=;/V9R:_/LXVHFLd6XF4PLR?JbHM,Xc)A+@
+7>SW@2D=@f<e<],.5>a\6DM7/:_?2<VMUYPIM7YA;Lb3)74A1F_3QcXRB_-6L6+
f#@N&?0NHUd&c&^T=,A.VT6JIP:f)g[V+UI/eH0D:21W^,OWaP0Jb&.6YLe>VKCb
_>V4OXPfIAI[ef-dG^4OHgBO#FMT@;T@31@Z4X+1-,H]A.aQU5/NY1FM?I;A1.dL
^J_[MKZXE=53gV/+gaIZVg+@K1Bb.DXT)@M5(50[g4G2[+1BF_NWMVIQ06]H_C,Q
bOaL@-Z.(HJXLQ1NS,M2,8BE-0(,2a]Q^+a:9&9[9MMW)48>U3)W4&S^[O&929Ae
8)87MS9F:F.+KACZYKe4Y1TODPR.I&OC^d&/fC6T=RS[(=&ZNd06.2da08FM3=<B
CEPa(+318:GKRX]c=<?F[Q(,Q+5]0^Yg==CI\JM/SeJ)cN5V3Q7_V25B9E]V9U/.
bcR]#4Y\fdK\^:=eg.J0\-Xc-EO_MfG)TVg,+06PG4^K8=[b8AX/KZVbC,M6P,G4
P<S::C.IYYB@&aE]a8-Q>V_ff@]S#d[A1DG8D&0;Qa-f(XE]Q@WD.5QbA]H82QT8
F(@=Q+7I9#JCIeaU[4Vga?:VMA0SZ404fP_/T0/7bPZ><TB@.V;;>7#5J[a3=/.>
_0?aDZgMK=RM3Q@D0=5/[?IbP^;3G9YST[0CTA#D;T/=KS:f+BU#W4IMU1I[&XW1
P>\c0eZHXP4BP2E.1F:a3[43/59fYAUJN57[&Q@K710Z5V4WBK9<Q,.Y..bW9LI3
MfC;b@M)ULZbIG^.^WJ0M6RSE;9-Ka?d20;V5G2]<\T9J@S5J(8/OOX0GLR+e^NA
?PcZ/@2U6gSMa-R7FAD]]d:>\[fIC3GIMGN(I_HYO?W5U&:4GYR@ECb.R=CQ83b\
d52#0UO)<,#2K+PFZEH&d]M<DV<fdcJ(ZI9:4A9UVcE76VYSF9O;42PL[X->+QZ8
O)NEW]S=1IB49#Kg=MTO=YH,H61UHISL=<eZ+b63SOC\LdZ<9]4B)YA)Eg66.J7(
OXJf8B:D3M+7<B:ee1Y8EUbeXg()G?::Jb_A@QQb[4I+MR+N8#G>?)S;eDS30Jgf
/UPecY6/f==35TgZIId59YQ5^EJW)@;F-a775gD9>X[6cI6LDA5a1G[0ET.TT4.O
<M:QN(GI52FC_7LcMPAK4RT@[)=E,c.MPKSR922ZR/=Tb\XU@SL]==B]YZ<9b0NL
2O]3d+CbQ61JKH@LN7;@?M\L8a++CP2c:GW7@AK8=7bfQS&[TfQF/EIPacbCBZgM
I3)&3/Dg=N7)I_c]1B8d.=T7Q7&N6McH;VZM?J):J-e>V9OBZ4WVbPG&I\G8#ZFS
@+CN,L#T0U(QG^R/A7ecK9_W^E6^3S82RXAaCHe:=Ad([1FT_718=N\4)P@C#.f7
dUZ^,(V6GV<KZ<BCUMN5G@O(#]5&6\6?cE.HO:]Z/LQ4C0&5>JK_+QJ[Hgf?+\H8
7&W?2QAIL(d:,CKcMA1bT.^X;?\^_R=6a\?7E<H+G[5W@)MS?R8)8Q7C-UdU@(9Q
<CPXaBUR+&+NHG91UK:2(IMT@9LfK10c(LcA?;DC29J4-72,?32LC[_eJTc@9O.a
ZVXXd\8F)?1R>SIV<g?[aFR8S^0IEQ]X5c_Qg\1QS5_)f;BaJCEK.Wgb62SHB3X.
;&ge?.0,A/@^G@/VK\YWVVQ[S-@K.caC-[V?1KXHWZKOO</b#^fa6JP.)U006?BT
X^=Za)+-:aGX;J/gcXYER,/XSGNL_7RWZF2M(GBA-S^S@H:@cI5>X/ad7XfMQMg]
PDT^gSc=84,cLGJ?Db@D\[Vb=DaJ,\,EIRK&SZJD].,TN,J[L.]_@]YgRbW+);:Y
<&VUYH[Cd</\QDaQ/]V4FAGS/<RB3H@^3gLfH-\MC6ZC:RY&(E>)1^#KJQ_24cbY
28,OY#>,O@<@]=I+W40J5M4SH-J[894C@TQ).TU]_5Rb4CaOg+6;3<C2.c&M,^P1
G?N6bLR]Y9.=6)5L4+da=<5C^FL9,&[2,O>\J&KEXe53W]cFB_]BW@5.J7JUDIY>
-0TU##e7CCQdc0W6.V9&bLc9?f0,6dZ>5<7G,Y3Y=NM#R#@2<8R7H:HNQ9a:^^ZU
@EC#>,?5(EZ2[[]FS0_]0b=R2C2/CL]:@S]V(QH8C;BKc(\UGNS9gV]?]Z3JTC[<
4U6OHT8/B]R@I)/RMC_IFgO#]?.(,)4WDbU,)c)]LeY@\^aIXG1O)QV#gMTBUMMY
>BN4]KaO0Ja^E;U04.Y2N4CM/eHe\:+-CZa[IF.MC).)RQA\ZDYUB(F7C2;Z1/,b
LYO0:IM(dcV3_-VC/-]A4EXA\4edVG+B_c<Z.1,FK;We6+>E\DAe2PYG,3:f[+(J
@V+6)g^c7@.We52S:9GJ+_F:FQOW[+&R@(GT(BOCa\KU0@KP@YeA<_K&_?X(1Q2&
a-=_@3SF/c+N7UK_L9ce4YbY/,6):&Q5?[E=Va<7QRNMb?Z4@)2g8&VFG46WS>77
DF(FZ],\6=4S=-<U/g3M7^4X0LaHPB,HQX?0=?M6=3G1>9d@._-?Cg2?4)]-?@<E
:5]CfXZ9g\cCQ0d;c217:dB[2Jd[^7@GEDR,S8F&^_<8>&ZXUFe(G)fHI\_22H<.
BA7_9_X?gL]10#;+;]F7ecY]30.S\,c):R8?ETB/BRNI/GUbLSF4>Fa5d.J4RDQ=
KTU4c9R2&E6,P3:2F(._+gED7XQ17[,)(.Q>F[H<YOeW\B7]^ZH??]7B01eN=P-K
K394JLgXT?TOI.<S/-8L2;.R9,f7/=&^L=gN>I65Y<19_(b+fOF,,N4298MgG/Q3
YO1-<\d0>:??]:U7H4C1EA#,b8>N:3K[J++&f[bQ42F@FGO9_9c[BE?6SW+@:T4Z
I[HgWCAAe(.T1DFbX8=;R7:D@]<Y6]6TT3)@.@5=)GF_2ad8VEcA8L8CZeQ]6?(L
-FO)D(3)A2:a),DJL;^^JNF1HbYD&TENPS^VXEW,\.M[6g#2(2JMB+9<[=C,KG=d
)]M<S#;1-bK=PHc&#A2SY>VWV[(f:[DQ0c.4TNY9:R:Y=EAJ&VQ/0?Ba\dAID1++
eQDLadAIg<8?C^31@K>D\8/CT8-C1/G.FN@(5VAbGK<_J&R3P.GVC1Q-Pe6-+1C3
9:bN>Q&.bG,6<S3:gZH]N\8R[T7M&3,Vd;f51/D1-V(HI3J2_NX;H9VK9#-U#3>T
eSaDW]LL<8&fG)S:Te3FBf_dS+,L)0,\3/Q+<Ve:<QR#,(W^D)?-d.?Td_CF<E=c
P)5PR@INP6M;+YW^D]WaT.AS<<Sa9)[BLTD/L)BGd[D],HCX.PA.3Y&P9RCD1aI<
<GO0BMfK@;OC0F6WFR0<+a4fFWHG.[F4=;NU.B#64+E6KV-6SXC:B;O;g,K4MG\d
9@):+HX47]#&4d;/#X+bLXcEU)(Q.:H&\X=]C(9+1cTWaR=]\+>f>30,9<]@6.3d
T46F/8#.?\M()1]K)b^J<6<B_K\@XI\)0\_L/dWP\?=08V)EY+0)Q.YNYVa?RBW/
(V@AF8(:M,_P3N)GH0.b^)d^b^U-A=_77Y2Sd7P.:(.0T;F>_&O(GFU;e9Xbb96Y
#AZGUQ+dbDHQcJ>&RS@#72P_(e4cFKH3]2Z--_Z-FC/V>=f13S)IL7?+@WU2Wcb#
FHE281JQ3^Jc;aPJO)2LERH=QE)&31[\O6b.SGA059KfNVg<AHZAfTaRgO)GT#J\
PCSgF#PZPPPK)S1a&bL5dV1[KIA-?MW8&ad^Jc26[.E)Kd1eP]AP1^<90Id@Z1B=
+g[@^(<gDg41UVHdO,+eBS2McN>MY_UW,/+[.QY(bCfWFB0ZCP(&3.UR\TM8.ZVI
)_[e^)NB3BM.&Q9F[PPM_7;=f5NUbaT/VA-a#_]gQ9K-T=;LDA92AYbg.:T4YQd]
AY_d_,/fEePAA:A,-)+(G#./&VU6WGAeY@4+fB\(65B#L&bB,#L<F-0.KY:J[/e0
1W3>;81e7bfP=,)IIQ@DZZFQ5AaBd1c&C+:PIPP4BZ-E1d5@8&[>?V,(?:?&[]M)
46B]=-WQ;@GVFR;K3,2e>/NCVO:O.SQWC_5Hd4I)/ZZ[@+fER2;K802/?][++bbO
]T&CTOJQe_L0a@.0]5-aWW=5?WQ6)W.]G@<JI9Cfe(VNXWIOfOYLGaM2M@=aR<=>
32,+5J-HL=\cWf8YX2LG3MG8U9W5&5CLP9H0?f.GDQ4Q+IL8_\X&R@7:9VE4)BZ0
JRZJf0HBQ2[&YEXBK0QY8KOJN+\U.ZeSP,:.bFA>/0O?ZU99e\TD8?7T[46U=2>>
)]PC4\=Da-&^D=6Q@1AbTJJ?W6&>GNfKV]WHfTYSD7g9B(9#>LfKf#b<1TOe?BH.
KL.YXLP2BHB#-EV1GD.5LQH=P70I/V^X;CVMY+XVT]1.GGW_/L#(U&D9OF?:O0/<
H4ZWZN:QAD:]JE0_F+O5Y8M1fOU0b.NLaBX.T(33I6eS2(aFGQO\[V^EWc(a/6NZ
>9,>Q]1g=O[.H\A<<D4_7]b#,;T>-AJBV;586dWT(&B40O26Qc39+A7KTPa9AYES
b;QVD[,.>Ga;WV./fJ3HN7Ke)+5fW\S]7B8a7+CK)>U3Da=EOUA:f9>T2P[4E0>=
?,&F23XH/Q&.UGg5]ZRH_SEY&F3NaY5GfPFEd1:ge85@R-#HBJ/Oc.A:+>&O&H=.
F0B9@acF;&-FQ;c[WU.S.4dE6,F_6&c&3e.SWLS;b\H/W/U58g8^_03g0N;5RK:(
-gHFI&Fe6NN(<D<P6bX6A:JBcg==4@G7_&XJ.a,SgWNJV/CR1O1c&B[aI^)CGO^6
J;WY#d-=DgO1^L?fS@UB)ZUF[aR1\P^5-,0>,_CR^VDXXRU#4Z//:@E5&@F<PGM9
_^(LdbO@TN9]<41ZVC[MPZ&C?G21YZPfSgcB)d4#Eb@8)9G/gdRM5g5ZJ1TRQHNT
KFPO43?0Oc7CIYXW0UZbR4L)2e5]cJ-3ULAbNJ^77>,bCE0g@aHV27;ZM(\SL.Vc
Q=b]9-<88fQL_S6W>UDTA7_-HR5H[Ee<F@UXX,\N?9#MH>bP2D&22Xb,eM<COcU/
CKZ\\b=D-Pc#RET;cB^MO@WR>6GS?EO<V4H-@JAP,G-d#X#S//\Md)0C,H,:fBIV
+Y(@1UC#0(5PZ2b=B/J\M4))=7A?PQA3#U8VYLf-P_bI-2gC=MaXVEe<bZJJE)Q_
-Ha[Vd(aU.QOcU@B)ZDXQK7Y[K(^]F\bP;bdfeKWF_FAfBXD6I_[A-O(?TeB0[B.
Q-E0E\Z[[N1)HS5V^d)Y._U\R:NT^V[Z<;\I8E]TZP(IPS,/V1GB)D^4A#K2E3cG
Sf_XL6f@156@SUHYI->d15>3?.^CZ4;&-+4K3Jf@GZ0[S1ZGTcbe5V0CQS&:9CO:
0_6]I&^?:#[8fU?e#A,R=]&@QCWO#eMM;Ef)D\F3CL<)FcHeH#c#.QKP,3+Z:TKO
V3A19Cc/YMQ6\4+2D@7g\EJ3KOTGERU:SB<7GVeTKcN73)Sd8IU#N@\?9>.a0S=Q
+YNTEZ;d^^F7IZaWP&eP2B6T83Q6X((-PK#F,HEf<7=:O(<3[eEG9\(4TC1aMQZC
Y25gU^b]6ee&BZ,=FNT_GLd.A4<caW6NBe/b8;UA8<7E#(J?BLLYb9J.0&#HC..L
d3,8?10MI+QPe5B:M_O4Qb/QU@)7>;eAO(T?,RJHMJdcY8O&0N<8eR]B7K[(U(Lf
c&PMU#SFGcc(0D?d8ZSDOg>C)2eHI)7E\1U9EKTKL21=O4gJG<DNL^<@,1APBM0C
;Z:DfD8#\Ab8\L9;;34^7?4Y.OWUF0)C:P3W6UW;-8F;;\Z-0,,aK(.4DOM=4@R(
QAM-?>X#9#(B?bH@R0)_Q02&U3=>b9G#8\G&(XgHP:5+ID0bR=HKg6>^^:(c\d9G
C[/T6I7N4OTZ)OS(NQY8(J[<d0f5;L(?7@YE64=J<O=360YeTd2B\+)1X+AGZSEY
[C2A]_66g8gJ5BIF_b,9#V?^CK:7B9FD2^Y&\B)Q6O&III=CB.OG\_2HR>4WV\\\
+:>35IF2AfY7P6NF#PbM/<+X:YU#6<XJU2_3X0#Q07931T<?24E/,]gX:/H_>6MB
HWIAZ8QID)e<89&9:1_RS=>SEbYgKO_.B@LD3F?=0g(/b80Xg.>JTJHR]2#DDIWD
2T;5Ve>RX)[WGU.]]Z_VBC#S:0DGX4Sa+#Y21OIV8+Vc;9/Nc_5MTM5LKHM.?POa
+M_E.b\H],4g?><<M>L;0CJKR9X3:N3MVTD[32&VL0\J\==b2FNEQB;HeE5^\03C
JUR-<eUf;K0&+fCCgO):>@)?9+-0&+Ub;^b.,3V]EbVY1S.-6O):b+a9JN6.fVTV
dc(fa;Wd.cC@TVGLUE19HZFL-FM@7aK6&#8PgIaa]fQcZL,E5^21Na(C<3ZMN1B_
Lf3FbTO;a4KDT[\T>->e;a=#0)B2+1G-M?8BKIC3O=W83NP/dT)Y^IU,ZZ+ZO#DZ
A8Q80\g5c\UEgZdXYdU@F4;>IaEV]:LR9YH#K#b)1:H)0BDX7f=eZR5aBU72+#=Y
U3UEG_Q+2SIaM\3N-@UIAAUf@Na2[3>Y9B6B^ZfU<P+MY<Y^HM/+NAO&;03LY=NM
@?e3b1>+4Y3,/E?ZOD\c=bMB/d9\.&.+2]6.YLeD68U]G-NDW]\2[aFE-G=?be\3
a=3\Ia+QP9CG)/U/U);Fac(>PdM)AbG52F.L0Y2b_E=CG2g6(L=RT7OX3a]3NP_[
@TU6F)Hc&EEH[\93:;)82.#.Fd;/ASa3M&8[@&N_ZPWR@,#Q._J[Pg[-WR@)56ZJ
TAS8WD59\Z&c)1\2\a@AM2KSU:^BSEFbXfBe;:;Ef<W8beR6;S4>R(gJ:48V3:Yc
I83#5..ZYP,BDNGYPIcQW84g&1;eTSQM#61R[V-LZgOPZeC?.[/>2?56bZ=>CU:3
MKe.HRK&8-.4@V0X[58V[J<)?E[9bd0;GO]E/@aX^dC^0.M?T+Vb;(ZKILA+3<Ub
&K&NfeP7G=FABO_PN<H:63KP#?eO><#@dFfK##cJgMM:#6:Nc).TAX82-C#BQ>;3
2-2;]FW_@HJ(</^?4HTCPS9?0])d+[\6PIJNHaT2XW8@F(M3eaZ<Nc/@HY.7:P:c
JE:[+W&UJ[<26=9g+E#AIB>X3<8_[<YO6S1_]._aCI_H\O-JT@Z\?-C<FNcH@=fZ
<<,b;OT93^,R:c.Q=GcOYM);e2KA6343=&3;EFG^6[6(d;JL;9IB.3+aS4ML/2T<
):5L:8V8GMC37MMUH:bCQc^)bKSZIE#20T4PXUCeM@8b\/aM.+L^,SPTb@NRT=-L
>0J.e[[g.b.]T,&W7F9/_5F4RQd_HF+UJb9WD;.H^D?#KN&ZIG1fGY>[AZ+gW]Q6
)FGDD<\9]bW<7D.>B:\e3D61S0,X=WO?bV64</@5EMd,_P[D^^&+7O41[?P5UQQN
;_2,I?#bZgX)42bRA^7U,]:[HTNPV2ReD7:g(2[:@DGAVE/>3Z/?D(\3W^dMQTH/
[<#cVPf8@eUX3IV.MV[U-I3aBO1VA46-+)U,XEIEGHa9>LTb[?/?A:T66J-=cWc6
-X^=&Y/>baY/UOPgZ:V8]>V;W9,LeV4TTX@?=7><]_1_&FPf=#V2ab,Q^[>b4d=&
V?Yc,VD<3@1L(5@<:FPK)#=d^g?C]0XLF:FbCK5]caYXEbHFZ9LQZ\@T@7S[;GF[
<:eK/10KG+0;2>f@=OG==6A9Ia1g@C<OYZXO[@MPX0;Q/)M71.99PG8T#NY8NKN?
eX0VcXd=@dAH^5BW,/d#81;d&VR3+)UII>F.,82:#U8:,Y[dR?6OOK]M:2@4(#N#
EEO:6fW\0:C6Fb4:D.C9A&#\(BUddJMJ8@E72)&eB_a@g&F3#H6(Ja+HFOg6c]@<
OC,V3?>d:[PccXDGS)D\]:QcOO3<-6447<f?<a&ae(A]/=b3ISbAFJZ-(1c[?00B
1XL,cOCK7Z:NQ0MB7Vf>]OF:Q,R/P\g+2-^4<XR=G1YS00RA2L<g/RX]A(FPD8FS
7c,3CLPRAKQH)9:aB/UT:O_]H+>M6+cE[T;?&7FdC,]D4_VI+F0Ic\O4Z)-fL2#J
GSWEW>I2#K]D39EcQJTCU3)D&g?)1AV=49dTLU>]WE+;fP5CKHMD\YI;=D&4F)H/
(X&22SQC9Bg[P5#EI&gW(OA:XV_3fP8F<4TU@1VJLKd[eZ2-XdS1:\\>b_EKNUJ5
G<#W_f2/gP7?/9=+C.KSHE=#[T[a2Cf9g]QfC4(Z-R-):E6]76\)&4Je:9QaEA5:
Tg-;?:5,KZ4;F\^(9HW4O@D(;L:?G_Y)cD8EZ9Kf2SF/c,e;bCW:W10SYW;(D595
==0)O>LZSTG,V;=7=Z-,LG7T(I:#?>FaU,+3HH[@HI9#TS<9g;c9^P:9Y@,Z5Id0
c\P9Q<BSHd>+QK-FEB[8>\U&WE98Z&8]6?1_O46c5+2G14Pd2G3^bf9YL-R7^f;M
3/-^G<8SV>\>M]]>)d@PX7_L=g/-c:3@K,W76BDVMM<69HZ[28?)/,8ZMJ.S6cA3
SPG@/9(:2b=LW+<G#/11^BTXH22K^?eT;+46J3?L^<VB+.H\:##Z<A5Q@44b))Yc
X^2OE&Z2N\^c#]3_?/SSZ7d<@YVf3T.TdQa1EcV?AB(f9]H-+T8<\)8\&X2):30@
0OcGbQ-Y0LcPe9U9]\NP&2;V[YZ,)S)3OR^SX5_8,R=,?JGEI(=>>ZE8]OH0,aa>
Q__E3UbRcH8S)BW[:&_2[(#[H/f7.gfW&g-;<KX)]B0E(L]UIdQHO]<Df6]aB72<
;42PBH?66+<)[<;>VT9(,3TPR+CA)HPRa\Y2;ADWHS_EN1X6WbZb47C8@C6BR5SD
<(,.[IL.6c?373,UN@3^P:9AUTP=8a@2RCf>5R6WN\\76FL\fU1Xbf>.51L^aQ6W
[<5gGZA]fH&FK67#dbP]c1I./)\2R-8Iaa6PAL85=/1WgXCI.LWJ:_O/Y@&6e\8)
>bJ=NZ64&/O(+cN<DeFNIS4?]JNYB01CdcTF:\T/E;(W9>Jdgc<U])&)/)9VCJC(
:,d.6T)7K19(00J^X_VV,Z2gR2ZV>ZE?^,RdeSG:c>a1B5/MVQ]EScJ83+2@T&CW
0>+U7,33Yfe<S:G[HZ:bT,VJ9#::JG@+Tc9V@cQ]V8Q6Je^8PN8C]G_A+dJE,Z.1
HG+#(4d,Jg0>B@SO1;G.F..XG,],SPK7V7KP27[bQV&d_0#T;P^GB(9f8+\>K;;R
e:\,S^<^^b2\SgH[+9MQUPTQWg&=Z/7YCWUU1H<FJ)3<]99.Oa@gdM\,SVJ^O:I/
Y2SQbV:94(XM6Z6E&JAPXL61Lg37:ca(65=&b-B0N4;8.[VJUX&9\[O=WA\VMaAE
KVU35SJ=21EN=CWGXNV+XP&e(T6YB?8]6/ROK-#-N\\&Q_W#6:AI<DI?0#()Y#?O
@^UK#7J7Oa#6NVKHe:N6HL9:TG]0;aNR=X=M5GQ@R74Z)fDeOB=ER+DJJbB,_FF&
RbIV@DJ3,[]TL+\D5IQTCI.LC,e7LZ7+4,QZDHUH+RG3ZP9H^SBRfO[]d2Ka9&e0
[4SA&f.<.AY#VcH0P^W\dR)X,>>B1EVAZ99#4CCCb4g)W8?M03+ZKNISXI_1TDI9
DOKQ;3Y(YXaH>_?68G0BF]gICZ9/)A]#,=+P<C&R8e^LO.8T_ZO2+T[c+OMB7f7D
K2EbbZQK,C@L\BQM&NI-Q84f5F(K,Y+U?dB>+),ALN[Yd7d2K7_Z>eGJfb#LC4EF
e#+#[MYg9=b(8fVcB&\^70=c&P]>cXPM^<B32[A.Q7;TGf]I^#XLa]5Q@I1=Z.af
:RG[TVVe;HM[&W4C1Xd(d3+H6TNKbM8#K&O;1[@0^)4UE.IO\>X8E_A1JR@G+a9]
05ZBV+(;#/RO]f.U_YIf(I=fJ7A/UF_[CXX9C.ZIM[4GO9[X,.FJ],/<[XKc7Q1\
O[&D@#bO8>;Z:()ZDS7.L3:_(d<V29JVVB;Z_gRHB>U_T1OR_)LYd-7MN@2Jeg]D
W#56cU.T5+.&_C]BP:K9HB_:PHMS]1)#ZSKWVB40U6OS(MXFX9<KNgGbG#KGc1@3
Z\+\&>3Na,G[fY/PC.2PQE3..4NM?_=<DdBO?R4WeLZc2P?AT;MXNS9X@1#Y@cW>
:,]J.K=9MA_3IFJ)D^=3,(>;.7fd&W6:+C_@EQ546?2HdK?\Ga_OC95BLXfQYYS9
:CX<]T:W]LB1AN1@/7R+a&3SR9e7Z=+0MgSEZ4ZcCB\TQF^(Eg=)244ba^T1Ag=B
HKFKR0.@9U64A2]7D0PK2]((f,G)>/Z-c=+Ga@O_Ca(,BJ,\/UI+IBdM;Z/>:&?5
(4^\Q2c=H@4S_&]8WQDXD47V<W8<d,aX]P)P;)c@<,?SFFMae5Cf15dG9NM9dDZc
(,XdO,Q(.Z,.23Hb7HO>=L-b6L+AdI,&L2YY:/-DR,21O0F+3Ja;D?W4:O294;RZ
<WX],KCfD;I_].Cc7ZbCG_M-<THM0/^/,(\RXFZ9/>dPRP7feD;I;AB]4OLG<\.R
Z&AS-BSW5DRKg.87(S@@&E@.@.8Z9D:8G&-g[fY2(c2L.+I0\ZA>1VGV_S>AQXXR
CbNXAMe[D@Ee=\)Q9ZPd=+fINB0\<JWEA8<I(AQXYeW]L26[73KS_g0J8^QACfU:
I[Gf:<N/4J\;FZ08YFP_Z_@(=<Zf(QE&g]#IU.b#C8(F]68Q]..IX=XIb9A4>O=6
>1-Tg#3AY=6b.=edK_U]+.D6dQb_]3/f1BTEZQQ:ac\A2A-+G2@3eB3/U2&cNZVb
\9,]TOZc1d-D@A[=>JNYIF8,TUAcbPbLEb:,&36fY)DR#]I[65RdV0?9c9;K>Q/C
XSJ@)4V85ZPY4Ugb4=7PV06K)Zb9Aaf;G/5(/4^^=NJSKT.d[gH:@RgJNcU#DJX?
O(>AP\g\Y8B,9PSdM_/,LDOKUdB.cDVcS0]e965W@63BWLYIV-@ULBHLC@>^fFgL
Ybc;5XH7TWO&JeZOU\C/28Z3J(8DAd.9&>9ZC2HG_Q6X5TaZ]#T&:@6+b=9GZBO7
gO&I@2UK@AQV,9DX(^>#MR53dX8EN(@8,(H-2dbY\e&f4STDXQ/5\<7<G\EKX^:.
bc>?I>-V?LAFHg=;?Cd.)<5dP7ZZQ31R_U=_3Q4/-OKVONR7Q-b0&X[S2B#AFQZC
KY,,0/8D_.>0Ge(Z_?,4A4/@UebI^.b9;35aC3I1KKPR[Gg)]aVf]2+Z1:JI(Y52
2cJ0YUS(67.gd^a^)[2,8f0T5?6KVYaP>3ZJI.)3\E[QLEQb[YT:GC>637+DfRYY
:C/8GF;@@.GDEAd8:11:aM+-@=eN^D[59JNG>0#E?<e#UIM#1/8]S\@6DG6K^D^P
]+V:+A.5?)N_fF2YL&<:QPH@?P.Y4IB,NUA5(]<33b_:7_K2HD=fR=0TJbg-gSc6
^a#M4g\Y?Ib/g+J3GK]-:09B^S.GBHGD0I>QU\<2U><=JJ@XKDa5IECdfH[QU4BG
OZ]_^PB<6GB]L&eLc;J,<2FRI&V3TQ8WW_^NKX5d7X+><Y)eRTO/HLNCW7F1b7L:
b9e7<Jb&cFN9AV7RQRB^a9WG8\+V8/?>bG&LV309#J:f=eJT](;T9MGRF82UfQ]a
#D].-#IYg;WX\aF&+e?cbYWW.#(_cH\G.P+VaX0DGcV)M&EHO1&f3W-T7^[RQ9bE
QSJWHKS+(+1B&LRECQ@S;)1^DM05D-Z-P)8C+TJ&FE>-,M7C9CeO0VJOH6fOUA2Z
eE8GZW@<dYK5H\]LYTRK8<-RZ_HHIaL#]?BS<9T<FRU.^?8-F05dH\?JRD[b+-K0
L6L:,+-5DV8HDF?)E3X2Z>CWYAC5b+3;J?B;GGR+0CJKN;/9F(E97\;^TD<7#G=0
.Z91M>F;M1=3@N9Zcb?/N9+JC(fPTYCA3Q.Z_F1dH\\/PB:[:7,-Cf+MRgKPV3K=
c+5J>_bQ,Ub?OBO-4UEf--<+KX]9);B>&P[2[K4dNQUUVdL4dPQJK/UAf]O5f_.[
GAf2BMB^8cF=D7U-H3HNFca2bf2#N],_.T>fH<;F[QQ)1=)fgH,a&Dbe?/7NUW+;
B]]eKK^4LG;Tf<T3(Q\3-[>1=P4T.LT7RX6NTH5:THZa@?g[0X<SKJD3CFL_MNbP
]e-bf7_Ea0gW._I^gfGN\D4@C4R=a?J-WQC/]B+]^3SW,H#P+4#9T(.2OH)JP_^R
AKb7;3&8&4OHFf3_=?Gb<f:5&9DUTYT+Ed.CeFe(T,F1-FB?JGYA64;XF/6@X+46
](KfB9/[)dO9ALfY.;^<LX>cBO]XCH<V69=\ID;UH/CV1]fceWY8T7JFK4ZIGeC(
.ZVVE/Ne+F@45dTDL473=MYe-2)Vc/&.b/RgIPJ8JQ:58NHR+b;UJEMgZb;];O#0
cW<_U6__OQ39B^MY>K96^27:J<S\&76aC_f-@AQZ@C3d48b?)f:&^NG;\92XHS.>
Y1BHFL-cKQXc59=74+YQD:-,.?U-C(P4=g1C4@OJeN3U>g-Q,ZBc55)=CKPX>3TM
CQER_JO3=YD.SBPC7BOC(e=]S==T=Gf7>HcMNX/S?P/?XRYSefc01S>Z9#.JI7YX
L#/4Q(^QWH#6DJE:E35T=Q;>aB(XT+FYUT3GIIRa53aV,2S&_?01HJRD]d3PKd3S
_5VCY^#FKT/E>bP,]N@TWeE7,PKSR=e+N<9<X,BM;.=,X.=RFC8C0/PJRaJLJ4gK
,BGd/#486eEBEZe.X[G>6;@ET[a9^6?UgX>(+g9<P3W2QJYO^cfCg1=U9GOZET\O
V0RPg.4c]YLFUOZd(5dGYR-]QU2O=@90/#cAC(>;AGN-CN#QL(UAG[b8:_#gFJ7D
cORBeH<J68_-Og\;eO1<KcY-D93K\&EO=Ta+39dWHf7NOUL5EJ[##A,RW+a2(Y[R
9.WJ;P+T4FNVg:--65-_ICIRGbJ=P(C-f17c/=<I&7FgQX)K0UaG>1AT)U[7N\5c
DWGDSH:U[bS(DbS,-5D/fO&Z95VCK[?4Fe755EMg?H(7XUJ^UH;g1?YQ0WQeKVa=
GT]P6RI7UfFb_XT8V1JCI3+)C+OT@BB(2.C.3Q>;2-32.G_[FCTNJ,/QTJHM8cFR
?50&3XSU@PMFEd?cER=:0\P3\FJRP\,<cT5N1;X<-L:0WfW^[8R:PIKNAc/aVZZg
AOa=0bU.?(fSZ-[P0I+cN1RF3g3-JW]cJ@=6+PgQEC;XF5^@9T8B&\0FWU08JOEM
.]2EH9L^\<4BQ(.2.P,Tg1R;UM)EVd<f3)OD-;&^&H2=d#2V[SX)5F,AY[\<&^PY
g2S0S.#66R#/D5NB+R?K-a2?aOU.;R.PK>D5B=^-XE4R52cd5c7Sf-F>>)P::5OZ
)9+N3>a/&&BLHOS05V9K)V&AE3?e.LL#_Z?5+DK_Kc]e^dLQJXI9R+MN+-#N/YeP
Jd,cfM_J.CXXb1DR=EV1,5gg2.MGG:(B0YWI=:\KMc6YC&4_KE3XQI?CI3BJ[JWZ
L9PDO.95.VD:X\++8TCa:2.]6Vg4P_O(X?7=bK;Sg[4;AK1O+/QGBJfJKQ]Z;[e6
N2QEMH;LJ)Bfacg_9-A9@?T><B.#Z>B+^K0[V)X@BN93OD,[[fV#FNEPfg^@:ZM9
A:N;:&)3A_>+U9Wd2:G+7I=-?P:,G<@9_GG5UF,/D\86BJ&A4PV5PFMcA69GR.-Y
gXI\5/.F9H<_<c1<5gJ)Ue2&?N8RIX-=>JMC#WNb90b(B_+c9X7&CdO=Ke7G>+7g
JRE..3[.Kd#?Y0DgP@(#;L]):YACOE>R?KfVHTdbD<A0\f7^KTDgd-cNDULXc0>7
ZYB\B>Z/^-AA(7M6[e_W5\=8&GE()gAYCDR(^b)+&&_50VVIV,AWDb1.;P_>-[R(
KZY.C-KgI9K]/WZWJ_<L\?YPb7b<<A:=2fS_7MR[8ULDT3/UB34VK[gFN@NL=5AN
TaTSA<W,acbf]CdaUgCNe#V;CY(E3CdFV5)093P5=1<[].J@If?;372L9&Q/X#:S
IHaO^0BS\TfG7C:L07=]&cVN/;:b,\3SfcKMX/c3#]>D@,JD;E3Mb-)M08ZO:T0d
5)V0XYW6[Le143e1F+?6/^V#1J#/CJC6eQU[g5AFU4D...TB/JZ,KH+LOgU=;J7_
^VLRWQ02]@Hg6_MZ)9HcGFV4aJZP(6LO<R9N<XSS_KFf1M>@)fdN2/6>B(YJJ4KK
aH.V[>ISK_8WZbdUdK7+AVWKb4/NBFaO>MQ>_239G9[=HfTE7IR2FIA32C^N#;A#
HD,38g=G&I_A+PcXUb]CEKZ>W=;YS(K<^V2W+T.]U;a:PcJK^OPY1R;@55Z3FDe(
7D+,BdcEY>Pcg?[57KGN;XY2SU1H)DL56KT/)R;-/8A<QB1Aae1Q3[c0[1NGQa?Q
7GVZ;OO=dQ6c@;NZ;;89e/L6Mc9_9Wg@TDLQGVME6@>KAX]RF@Zb4HceTO7#Q0(M
cSgB6Cf\WaXbf23/@M()8dG5U&7bV44MV-G1_>ELWXC,g0+LfF#-9E#RUbdaK)cg
aJCdaBK<,(D1;4#XBH8K<^OCK^X8)915Z)Y7/Wb0I61Z59G]fPKO=&ZS)f>#&\SD
bG]d3=.7Ob^07WF7=8ZE:&b9e2fD];:e]eP_@&6FgQRK]PNZOPHd)_g(@QOd\PJ1
1f>4\1THeK#VIV^7eaH2E#S03(\O?eG(Y[91V2J:]1VI^@5b6418QL5IUGL[d>GM
2YPW+0f&?F)7FbR(1C45(W^YB91P?MKFaBXe-K7g76+bMF>VAGH8Te,\521fCI6;
)ZCS9TDfFS3D\_L;/_112^;Q-_1LLUL#[^G(Ybg&(_:]bgV7HX+7\Qc;I9HB^I]&
QeJ^7C>MUD6e2APd@O?IaU4/D9/3,O3U,HT>EKCZ&.??[LX&CDf+RIaL>U_Q-PQC
,E;7)4F5JO+DQ[]^Y#.b(/HG65D-3&PgG;/VXZX]g_]YbUEb</+&:fN83O+HT.5U
PW=[^J1@J)Z#ICLe+=3STN+g:Ld@RUQd<K,US<^3Q5]C3d8f5^.-3Q,AXW\eC)).
.(RRMN\&>U4]e+Ia2/d(TYX,E[U\JI#9HYKTI_Ga4]J\Gd&/_@&E1(P.[YdbHW^N
G?.YZ_CUVcG^6Bbc(O#(X^)6c@E^0^R_b01\WU4]/LU84a8=7g81aF]3c\TXMQcf
aQ58/,1U=^BC[<J\9M_/6<,5S#<M&7VdUKCV(\1OZ?V?:bdGSQ1OfH#T7ERZZG(d
C.BWE?<be(35N9?EGgKR]ePS-,QJIF]7,(cN)5c;KAd146?X\\g_B)Vf)EAbfC<&
TQYCJ,RZg/gGWA:e3g-.KH3+^O+CFX&:M/>(#N92WOJ=,/B+eP=R8HCF]eI]8]U7
1Qg4/L8T,<JIN,AT><g2e6Z6/^Cd2DZe/CE=PE9+EXYcVe1U4D)@D7[1(QNSTHT0
,e9NE81SB:N@&&JU8A-8e6HRPROTC2T^H<dE02XKcIFe&>VYR5G?:D_OD4Z4MfaM
b+@KLc_<-F5SP-\./1JQIg>47&;.:@X-=]7e&fL3Q>Z#?Z&AR5&7Q)_98N#F9V>H
MZF-TUTUJV9g:T-b&K;K7RP3/4EX[ae&:J=[8^^I-e_5G13bAULA.<&W79?RK7IX
?e;3K[8UYZ2[)bc)Wd2g9Z(/BPRd9/CE30DWbV9cgNSadO2(8Z0:3b>-NA7F<PD^
dgA_9Xd>9-cQOBe^](ZcX3(?)#_?@5TJT&O5g(S^<AKb_bBH0&U<^R#GT[\5X__:
;CAZEEcMTWX#ACV9^YG9\dDN0(QRDRM?NK:SU-cK/cb1,Bbb@SY3e\0.0T=OI@^1
3IYEN>aQDNWIQ.).XPEVa;W?U8F&FRQMUUWgO[G2?c1V[KKL9DZZYJQEH7AWEB+-
SUJ6^,6][8:K@@,4ZbNgL4VN-7E,C(+.&&O3]^8-_EY-C7MP.EK=:e.<0;<I]T3.
a.;:@dUU[#@B-1CU_0/N2cNI4/+EJFWJDF;W#?QSSU_#IVH+;X]8_-(O#+a[K;Ub
^)[#]f=5;Z1[\3gaT9RM5),J<Recc,X)JV)e+Mc8=8b5P/2/ZVTI&4=3[25N_gL>
C-N?=#>E&TdO5H5^eHb\11g<[FgY952WGC<-Y<A8)O9c]?UT:P5+e\347X7B<3-9
1,6H(7O(OQT/d:CZ1?;)_:01bRb\7.I0=8R^FI/BL3DcHDHL\]/5:+3X-M9K5gB&
@9N_Jg^.BV1d_DQYg_,O81SF\2_>P+?TWMeZD<K9FbOYYdQ.4>9/P;_(MQM3RI4E
MF6OeBG?K\-C3V(_^QMG\Y#]Z)=HW:M?E@1J?B<4SDM68Cb4R+3:\W^Sgg6.)&Z+
Ta[.W>P#9C;]\HYR+>.5B>UY?NgO?63335I(:JND)_A+BB=Z=T+M;@+Bd])c2EP2
S\744RMeEI4;]1FQb&EMVU/J^-_3^2]YS>]MW2Ya)[D(TZ4H,+2+/+1J+61O/.;b
cO6fGL/EWW26STgLC3N9HEKAD4c26KPHIH.C8X@JCC4/Y-_<eIV-=-5Y5CX8+1+e
ZB4MOcXZ^12_0dTeAN8+TO1HAK;VJcMSJ_@#U;#Ref6YEc7@I2Q&e@C_41>&0M[I
/H.Gc?;KY3DV-G-C87C>[,37&F55CS_(S71VI1a1E;2Scc1&\fNFIeV7=fKLK@_M
J4Bb#Ka1+a/3-9+T1(E@[RMU/]M<M/C:/U9MQ:e7G7G@6F?H13:8d)I,\N([.=,N
I?3_P7]f272:#DK>D;W6/c2@0P?KH&9Y:CF:L+S.Wg.F&-RAP[&-:,LMXM<GN=\U
PR[;+CZ;@^V7X[+0O6bd2Pe[UOOM.[]JaDcfM34QFMaM9O\4)_[S0&O3UQSg8<0E
)J#3MSA^RM^NS-dAgg]I1CIINX0TK8:[,L-\[=;@1J#L[?Uc3/=>[(g1/N-B_gI]
K@XI,2I4Y/D,5[3H6O[RBf0?P<4\E=XAJ:cO8NJZZg1>_AUO(]&==WMA=+QXWZDT
5;(P+NCgX7XBSWY7gXI\HYWK3bY.PRTG6D9C..4E(Y&5,Z60E_D;_ZR03EY_dH8F
EUdHU^HQ^=Mc.KALZ;;T04)LaS=Q;?[;V_F?(H/[C&>&-OUBD4\F>dV+S-5F],;>
UfX>;Ge&d6&^;#,dUQP^N3841@+S>:=TB=80Y&\K^R>#&YO]^A)L)EJ>Y=R-M0_5
f[f6AG^E>PLV)XAN.Qe>D-M>2PfF[8.#/E;59cAZ8T.B2f)d-D_Z9d_]PKf\8-(0
.YXD5bTeY2^M])ACGT6_0@2c-YYg<+-5-6BO,U;J)#\6gYB)3\aM__L=-OG?1WOL
8IY=;eL?&/Z]SG:J<GSO,/2(14S??_P934F?<;g0MN\D9eDb;S0eX#.53bTI76]F
[BfAYEfC#;=\7,?&d+-P([PHAcQb+eggb=>W[^&DNfWF#B-3f)1Y7He7VX>;fSYX
C\Lf1J5\2gd^+X6AQRg[9af8WA@>1.D\??]22-La<b2_ARRGWH>#g_UgO1QA_4W+
]Rc4fVM@,M9+L#BX2S0b+<\GNXb6\[7=NI5?R#:]E]AEC)&;7[Z5U83Bc(Uf&d=W
.=V@L-ZXc/L>#OY-?_a(?-,)>MYJ<GH4_D\+JMa:^XE2]2c<2V(7b:XQOF)\(P0#
9=Y7&M=eRSb7J8JGLYQW)\-QFLTV).FJ^R;:@\#(+@@J,Gda=_]C@Tc)UcEOaMO=
8+7dU:WK[&FEXV;_+90[Yda;UA7bHYYHL?5-UD4G(I&OH@G>VPA:EC>6ELM/&.Bg
.<H;1b1;\,<e3]6cUaeDJK=Pc59F?E238R\8MSgKc:6M;@3D-5W4?,;CZEGM#3N^
f<#d8\29#\X0->IfLDV32cR6;Z>C.3eL3fQa.0CPK4JZ@U\,[Cd,(g@Q0SgF^2_a
-JY^0SI_XCX0^a80DMJ\+-R[SQfFPE\5fZgPR&F(P.e>@0^cg[QTJ_OCHUf/H^C>
)8X\]IS:[AC4O6WB1EI5\YcVUS-9M_O7\#3DBP7#4T2@HJCRc1K7OF[<7CE&73Xc
@AIXDd5bK.8_4I4E?P4)D>K&FJEe#f+dH?I+H#LE\/_WHR<WKGXQ?Q0IGR)1_bVF
83cK(N<A9#Zc[;/0WbGZ6b(LF0DH5J5?MHE;>cAQRYg3>TB]5g-3Y_>9SNLRY_<O
YQIMC8B?X10/?3AHf_.f,LP]PBG)@dF^_NBK,faH\eO&aAH<ZSUSbQf,1S:^GSc\
?5O:9L6B^>9f44YcaB+EBM[3ab;WC<fCb-^/6YV,^:I3J6LMN)#VT13R)4Yd=3C8
37A9Lg2R/E[g=?&b>A^O-^1^ODD^3M_0R(K^3dO1I(Y.N<N-)F[<=XKN6_0dUcZG
GRE]):U#7<S60+>4c422=H4e#5fN7,CU9E.\6ETIP9XEUOS#FV6^+P-_3DF18(_A
L>Z9H5M]b7X#1#U<MSSQgfW_(>]#fYS9,NT2:G4YH=T<PBf)M1@#B#?:fYXW.(SN
SNC,[,#,DS]+_F;fA7,+9@QL?+N@.E?S8/6f]H(^:a7RG8=e_b5N.YT;B<;?QZLK
([/IM=FYB&M0LA3c3E7BbKQS1Yd=bAUE>1K[E\]6W^RPgS;7ND^d,Y;HZQI;&)b1
[8LRBVa(7cFS3#(ZOC7G-fe(I+bYKM0Ve.T@AA3&ST3^/WRI+OTa+&a3BEIAK;aV
,RQbGOHVQ>=KGW8:76)TUO\KQ[>:Va?OT_\OW@@ag:]:eTSTT@gA^GX0V\U9J\T7
e],=4F)D^5CTL,#@5-?BQg,NR^X2-AEX?YX;R9B;,)-cF1F2)S/5\Z-fTAQL0YB\
f&&+f5-:WT2\DJZVI5#0BUD/55f,52C<4CER;0fM6/07J@;R-C7NQW+&?d@OZW>f
P(9XUeL4cYbCM=S[<ERQ<Z8_I\Z,VY:&IM(a_WGd:,bB+N&>;5Cc,?J2^)be_,KB
EW7XaZ:ONI]N0aJJcg/OI?^L1_GP\5U<>4DcA)L.?GC]Tg/D>H.Yg2YX:IRKa_Q1
8[I-5U.]3WA^3GJK[&A&QcV^G#g,?bV7R1QV-Hg:C[b+Q;/a=L\Yd3\;#L2:A/c2
W/)L[&L6-,aOKH;(_d\[8dPCgAY+KHGYS5c/6Hdab;_67O1:+#0A8=+(QH<B(KSG
G1)cM>XI6B[)15[d+G8Q0Q8C;(e&>#XX?Jd@SV_2QJIbAV(,af.Z^Of<FCM[8IO4
UMB0(;X=-A/TS#4=(ED+;,>cK0Z_S;]T[/VW,HJUcQR;A2Z:/Q4Q]2EL1O8-61<:
fEUV(4PB31_b?UT-7:0?A8aT\4#c9d@@.;bN<QG[)D+2-g[dJTdKcVB=>-RM\B33
>?:(U6.ZDcgMNI#S/8H2H6e;;cD=Z+XTOIN]\B2N69g=TGdXK1g&,Id0VX@9+c,Q
<DJ\aI/642+L>0;;6Wa+_^ceLGGZD+WgZ,/5=LWYFB.cV1VK_K7C>W?fT5ITFC8^
K-.3G3_?JbSGUX<5dZ7[F&cW\9TTW=T04/5S+E5ZZ?M[8EYMH62(f[NH-A-.KL2f
WXCBdO_=a1@c[];ID0Q0F(E:63/ND4==L>O.Cd\4RY)/V=K,RXI<9JLQaP63I36I
/1+.]+Pg<8dca>7>IU\cZX\>9B+_#N#6(5RX,gKQeAU]N0?2[C6;eLQO>8P9MJS_
ZG#EP27fYFAOFN-OUT:5_8YX(((.Ff/d5cdMOYa<>a(:\d79O8I+QaI&B)O(020B
+I=Mb,+PGAfHD[[B&R4+ePb#]B)^RJVe@(Z8T5]VYA(4Rg3IeI#bdLJVZ.4-[5\a
&E@C9:UGa,[FSgWS;AX9C9?DI[2BR-f<^gXGF,U<10S[^GRIN,[J[=#G_aI(a.G1
1\7H?:+B\#;U(0=;1,C=I6YPJK0WEP@E[J1b^/I58XJ>J.G4KfK>O5&J8L7E8@;f
;<ga-B#,2-D2=[&#_)2,AD2Q_-2cfKN3[5F+.B((-8bGH>])O(g0Z;/5^(b>f&NW
gcCJNfS52)(&MUb4N[]+7W8@@V>J7BTG1\EIVBf_?e_5:EL=gX,>GN1Ig[S1XIY/
Y7^/_17NQXA;YN:/;9aDCT-8d9H2I?)78>2S\_QG->F6MR\+SRdZ=[.>DL.N+I8&
1,S)fgK6SKWc\P8O&?81]9Yc3MPdJ[4]_(KbX<)BVPb8#JBRgHfRNe=[)DPFITCg
f50Wg&RAOHGSE^Z.:<gM=/VSb10=XE+=UQAM_YaLEBFEcSY(;5^-VJM#T08V+(J]
&B=#5Q3_8#^8=Q[80aJ.KF.)[=&g39bYaICYUWD^06=.P#<S0T]/URAD&94FJZ[C
]dC[TXL@X>MWHYB[-;E,N:0XYO1PPaH55I.a2+UHY3>0OHZYRbJE[#a?(fF&,REc
,[_]YX8cD\>f^ePB;a0IMZF&RL.IOY?f>M]8CNg56BCI_+Fg/g4R,IV-YPDXg2:K
J692]V8J:F@D@3Ad,fJ?N+5V>Vd(VaX)2c#dEQe,\fR9=&J:_2(D0U5d[RdACTMH
@@S,S_F6Og2Q&EDBZc;0^II4c)RbE3?\:&LXQ,SX4#?XMQ^/T8b<]E(2K=cTFde0
fHH<K]^,5@LR^aVUM);B)3EN>TY^f)0dg<d/H&:E+CZM3>:QJb1Q2GVB/@\:b:>,
M902=@\1e.g3_9.DaR8W7=\T)@KHBFR:DgbABPKIQDLPE/U7b>)JV(Y;Sc,E&(/B
;TO:MX-+<^S,SVEWQEQM@V9(<@4BP\[Y<J53XGL0gA5J1Z3>Mg+L,O<H7^EdXFP0
\I]KEJ1agBI1X3gCDUPW,,beUB4.Ueg#EEB?-3_FVRCWWM9)EXFEESQ\4@?MOS>9
7FPA6KL#+7)SL##@RfVe]4e;d24dX[B6(<4Vg=8U<1bFHBc8GZRLOBQZ[aLUgH^J
e4bH(<N2A:,X2A=-M989^RdcVe7)3/>:H1&a^]eWGD].L8D3R[X<Ie2O:I:7@.#B
0JWaJMC^P>C-Cc,@0D/##dBBVYCI4<T11Y#ZC5E7bIT=OHe?GS]Na6B?#?[<X7G4
<IdUX;]bHOdQ2:9+Ab?,&TQD9M_+J^KA_@+/BB9bOH3MSV)bSP.S24@e]G4Sa#a8
/fQ5:AJ350+\-5NGGWDQY+-++7),8M85K\R#K700IAZ\M0+S3].O-K)&/]gDFM.>
.C_]/a6TC](WLf#P?bfM;##6<KN=0^21Gc]N&fGJdNXO9E)W[HWS(MRW+,#&VHe?
=15W/;9\53245T;R.U4N<50+(=O1MO/Q7dG_Z3^DF+)LO38;bL,af9XfN&@#7Za5
4CD,16&.a2A)69cE./PD_J,J1gdZV;Sb]cX/7G#PQ.7,M2YHNe2UM7^T=W?@_1.U
H-B:F&80[<9MI)0A+F9=1\c/=C(,JW>Ydb-K0V4aJU?.c/X(BBRM=&4O_e]78N/M
1.H<=@K-8F.MU:MPg@M1b31g];)(98RBA/eQZ/C),ga[6]IGY/Y]bGeA6\3=\C/H
b]5>A&:;HW76@BaeUf@.)c6?&05^d5--WETc>eV,3MdG]IH(/DId=eAO<O#AaY=M
+9=U#UZ)>67N,IV@<J)#W[Y<^;GT:7H0_1=/6/9[C8XcYSZTD?/TbFFL8c4-S55[
]YDB@#e&<G9QLX,+]RLGUN]71^G@:R6\(UV[^;>gT&0VcR\Qgcf@=WO^8I-ddT<\
<gFLPN)BXbg3G30])D>U.gT.FX.X14R0]C]1\.:a[,NgBOF7bVOHOOb4,0JF[#/(
,DH>:aPR:ZPX\V9Nf=I?LP7MdX]0Gc/4TI#N_RRRCdFTKY@g_ZeU7CaFYD(X,\WE
V[ON#X\)DPJTa>G.[UKK0XN[+5Q3LVaDc9>ORCG6A990X&@K.:?Y/XBTG8V136,Y
]D#JB;.[Z[cebG5VN2-&>2XV[]39+IgMAMAbc99:C<defcGaRH;,NQb(@7RObGW&
XH[VMfg.JX^)FIVUPQ4QG^D1G7W->SB_UEEc\bQ]=;)MG21?1fAV-GSL]<fRT1gZ
GD+^C<fLF0?ILG0/\P)f=5A@.+Cg23Sfag-<U=,]\I76f+W-92P)gO_8ZUPFf51\
c8F=8M<L-,A-gZc2TW6M6Y&62N[3SQKK5+#0H.Q-H223D3d[M&9(;)Eb5dGF&S/-
>6:-581^R2PX<gVYUWSDDe5d&<5Sf>MK/,)J-RZWeF=6=_[L8UQL7e_W+SZW527P
EUN[,4,[;M>+=]fKM0TaN;7C[eBgA3PT8TT+R1].UKNLD3CdO@#_0ZW44O:^X>AU
N[<8VZ8W-P,J?_1fD]T0>;eA@:SLNIb<2ZX/ba2@ORM99<R^L]L1#b5HKOODBBE4
a9@9<N-+T\bG:ScX[RX;R++5(&)ZXT&CT:&A^[05eM[6X6Y(7T1cg[1.f\?1R7<T
BO3A?9N2AGRF>K5CXVED>)9:R\\YKJQ=;=M/TKgfRIa0]HVUdPXLWJ6V()7&#_@F
,@0bSc(>Ce^BZ:FV+^UPeS/;?g+MXN3YG-.A1VD1N-+Y:H(14M7TVH:)XXSR=ONZ
&3+4\3@f9A^;R_AeN/Ia]_VDdR+#TfGKT)_c6G=33F306X03Xc;;5DR,XeXX^b:^
;?T0[NI=K\F:VTPXQ76LM&I02a,R3.WZ7AbJTWR26X4aIJU_P<e;6PHJVbfAYPK+
VWRI]CY?UU0Y5[7].Q1O]&68#=FGB6?HFI>#0REM]-K7cZ?3Z8T;bJ,K-bI_[2V\
1_T(f5L.,]A^87CB_W3W]g:([>F=VX7(G(T0@_GcO:+&7c2^A+9F7T(PTNVZ#e42
H@CY9127GH>WWJ2:;ROW@cd./=KTYN_5]M(LF/7E40PEJXL>V0eeg;]OL104eU[4
D&(O+W.J2cLeS614,_f7=+K&6AP7X(<2d>9MeZBH2O;8a#WfK[eES),T_?b]1GUA
Cgd^Ab](#gT<MB_P/;&;f<a;-I2&MV_17,_UW1AFfG,5<YB().0YbHCIWXaBaT5A
&g;fC4+<_LZ;>gg,9KCRb:HfV69f<9Y8M]J,QY/5<&#+Z+\9XZE9fe88UE/IWZKc
\PYZWSU14SOU=[GObOc8Z8SD)4I&Wa9e&+PEO8Ia7Ga@ef7+SN;DQSI/eW8OMX?G
<,B+NYL\,Wbb5I8>VF]K+/=EAEQ=bI=OQ9gR-NEMA?BSCVDN\;4<-J]\,[E3U7#d
\3E@:9&4M/RB]YV#LSb,30MV/3(@MXXJdSF6_0FAYfW4R1.8+d&V8IH=O3OI-/SC
G>:]AN]P<>W9(#I,XKd+&HJ9CDB>)F6XV9V=c>0N^?F36E-#4\LR\E;Q=][1f/fB
+Bbb&XM.(T(H:.64#fZQH]dbHF:W88G8@/VCH8V.+9,PT\R:N#cL_I,@XCX.fOb/
DMcf#/)18S(NZ/ZbIb71-/0MM@2&EcC@D5?Q24?>aEeCD-3>,7SQT+<\V@UXI?<7
_6ODSEXJMZ7cV-5ZfEP-7\/0US/=(cK582^Ma]0+-CIgOMRbZ5.b72+#c?UeM9[1
#4]20>Q_Z@/Vd/4]3^a]=K#AZg]_<=ET:KNPa7TT1L1=L,f+.+R,J^>5-#LJ)Fc;
W9[aDbA:XZW\9XU:D,9>OC((3@[b\W1\YDW)S&Da5;b8<MFL5e>KMC2((A6^JRI-
+JV>b:GOZHKO4A[^S)-2.7,U@3:LN<]OJI>DT&45/=Ve=(M08UO[)a?+E-PJD>+F
cQ)A0VM4H47LH7U3N@Uf]>_S+&U.BC^NPGNCS]1B1e,VD^TO&2^DW&409-;F67J^
7_Y8d_[8K,,fSb867:L?/O^gXL65U,#+(BG;KdQId;CTF1KV1U9DBe8>W1V.KW-Z
CI0B8be2GN9aVC&b0QF7fDJ7^T@#eWa<b(FB2]@PKUQ9DOYHe;3XH5OLB,b,?(/c
Xg3]B6NH2HO,Sb4[1XfBYdB+2_KKdCdESJaV?CA<4FC/[CC/BFBcH^.20H&?eJ5b
)GM/&E1]4Z=],-3JSJKf2<2e,WSHb#_(XTVF(JH;IB>Gg0;:P>G\g]:M7R,If)\f
N#(J[RQeQ-#fJHR3])IN#D=:1#F)YNAV1.S[\c##TF?CZ6<IT837?M;Z=JcccR;Q
cK8<a[HO3Q[##MJ]P(JIM6I?+SCJ/^cN<WNS-L]&SC,/DS0GP@:8fMNODJeM4]2=
^#A_1T?KWNSPL5P8B[ZYK^e^M)]Of.6P4J,/>-eKe==0O2?^Yg)Lbf_<MQ/P?LS;
dLELWbZ^/<NPRM?6?.]g;B:I[4&F@?[\f#W<fJFCF:[@-]S&K(0D-T.0R8+e-O95
#UdDT=]V#24I_-8g]H:K,#+@Q43ZZa1_RR:d2S&Y:#Y>OaMgC+<_DS0M4gaJ)GfI
c/BBUJ0=_c=e=-fIf.UA,\SK)(bbV7.]S9cKG08X5@7RLRGB;e:N<QZ6FII\,2Ua
:57b4(3]3R>OK&W(=>0X;GW;_H(PW+]C2+VI93NQQdI]Z_AR7PXE.)9I?L3[V2A6
__&4PDY=.,aVHC@=-M]-ZQ4?F/e]K;.C>QA<8@;O6)207E]#=_PRW>SbeHFV@QTD
71C8g@XE.V;S+\c=7P,2eB1@+c+^Z-dNLGV-CO;@Xf/40V[V<+,FfPRKHE@cDQKZ
>09IcI,fGa-[=\@f&O=+8]JG=RZT9=)Q-/N7_c_YQZcI8<S^D\071M-SY269bbf6
20VN7MP.OCSL;E;RR_RNb56O/+V?[@NcK>O9GNgEY-8dag6T_FZ-RP7WZM,H:M7^
9C?8UA,2.5-[_4)d5#HZ:@R-9;C:VYWBDZ)47]F3JTdP^<4gHL9:e1LN)U1/[@a;
7V>YF_:./[5438V9^c\HZY#GI882O90H?)DEB.AVE&_91f:VYO.7J8fHY&FL39^2
+GC:6:&);B=LcXU3FL-O@_:G)dLL_&R_NYH,4>Q4Cd/WMgWgcC)DA,OXSb7+>N6H
:W<CbQ9&@67;XC(S\:V)aN6&52P,/ISTf<9Ieb0WVDTO7;@,T&d6,\S:Lf#Q1M[1
P@LEb]_D)@2L;\JT+7aEd2BD?6Xfd/d#EVI\)1-XQ)-GHAZd?Ha;)Ug[UF<J^dI2
A#6,<T#cdX@K.F+:86<G6W#B\P=PfZTc35U+3e8E0b++aU;AA=E7F2>\G@g]WYDW
IZ+II5;KTH+V?T[G3cTa:@e3H531W>L5-1O6=@UV2II3aH2+\1T.QQ7\G.TXQQMK
SCf0X,=8LH=\?g\1KedB2QCETc2V=D7LEF\Te?7R<U4IV?bU?;_X-,bSB=R]YD;U
b+41LYXWN_dL/?a-=K/?4(Z04/.M6MB:V4eA;+9?C>8XZNUX7-a@XFC)>&PLCa7V
U9e3aUMO11e(LO:,5X8.VaTTK5M>G6&\9[gBdX<1V/)UYSd0H)><YM.^0@SXc-BN
^aRZ#F\7V0d_</=R)=PM&8]<&I4JM?/?a#0Z0C#8BLJaB^V(J]?(4SJPB2E145J@
V</-dW<1FCc&M&70OWL@4;>YRFV\K(P]Z>2[P_C(<e2cI8YF<J(&>3Q^1YZQ8O,T
VMX^PDFK[;C\?-<a)AbGFZcT;VJe:.?FYIBT97U,Q,R]V5B;>(IS[O<])]dF4a^U
M0&FD7a\a56ADK=P1:4Y:ICR5NFO>OHGPS8#T[?>6EZ+[1G+EU2UMLb:LZg^MUEN
BH[d@f)QTEOJ9W<ZXK]83<fbF9Zb.#9W12cPg;;/gcF/L2+fcTV4c/,HdO3[W?KO
2RXWG&+Y,9Zb]?-Q/b<TN0FA>#F:fW&]B^RB&M>@FKZNJSL2TK/&L5MTY,0BI/d3
[b&/&[KaH-KI[eEJc)M_GD-N)^C_[)6DZ>db[IVOJ8IMOWMHV-,Y?d3/UW+#_:Ka
S2b,(DJ7[^d8->DeS?)T;geL&Zf)OdPN.99g1QdS,B-Bd/B9Sf;MS1d&9NI5_;gC
S0@+NPX/33F)W[Y4)1K7ZC@dbTAP/Z_.b@#T+Q&-H7-RE<N]YN&bE6SeWW//V3NJ
LZ1828:G(3f&0Ie1aJM@?/TBc\LIf+W4X&0ZV8F._RcAc4#PI8GT[QQ:=fc[[DI0
K30L_=F?(,(ZB\BcZd(TQD[/RWBVW+_.JWDHA.+1?\QfE+A4X3\.AP)O,??/;F?A
.?91^_.ISAJ+6M5Cg2gI\a4#E\WV+fTF&M,>.@ZaQ5Vf[_3:0a^\QL&+GY^3ORQ_
A37531Fa_f\)/dKFaJ]UE_I-C624\Rb]Z;R+AL<K?NL1#.VRd?C+:a4#D3=DTD75
W<VCPUM2\@aQ.V&V+X[?7g-7W+3KMYf:2AdbLNMfaHc6169]d=W)U?eT<3a<bK5<
8e<]DS?GCDV)>\B,:EeY#TR+K[I_ZPWM282WO,;=76@043G:4c9Eb2];R+147)X6
W#fMR#X6f#a36E/-:2/dU@1^+ZW+P<]:SKfFV_@G,2U?d5cdQff2_M,eW+B_RdV0
Z3TD(1MaA&/Y/O8e&;EFZ&DL3WR,IA@?07-^4:\K/E[&UR_90X0b.PT5WDBD,]:S
F+:K]UcgJe7Z^<=X-DGA:]H-B2Z(_8R+@6&KZ.)eSMH&A$
`endprotected
