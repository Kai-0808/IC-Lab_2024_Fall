`define CYCLE_TIME 15.0
`define SEED_NUMBER 19385032
`define PATTERN_NUMBER 10000
`define DEBUG_MODE 1

`include "Usertype.sv"

program automatic PATTERN(input clk, INF.PATTERN inf);

`protected
CO7ce9H?1)BD/ZHIS29E^IXZ2NP+.5F&GD7LIIa?Jb2.IFA-)VF^7)C[V7M,eS/\
bHVWG&U(g;(J(76OQ/&/JCcf,59Jd^[PHQ(RN-K&GLDA<;0LJ>K42,PK\U/M68&8
H9Z<8A_SVF##_BBYfGW)7?0@>(LSPHcb3Sa\.J0g>Xg>=65TYKIIK;<LN+W@;_dG
AIY/W>G;gAWA]USQYH@M:B<N@=XJWR/(+cO.<d#\Kff=g8e,4XL()#UFcYcHKENf
Zba]fCS0Bg+:(0Z:1^[S&M+7U>6]S_d^5aL6#NW-eQ68KU(X\#c27PC,OaHg6A-d
X-RQ>4B[Xa,2[eYI7AHaI?(2U<)72\1b_,#3d>(J<(Xae)D0@5XB<?4DS>:L5JWf
Q+H<7CQT1.QIY3,U.U?b=;07])Xd3=^ZVD\T\OVVb5e-]RBKP(B3S6+4eS+aaWaA
HbTE/>Z,gbXQc-c\g7;g<V-&JJP:DCCSB7^^/5X]:K6VS?6a58Q9PT,+eN-7H^a@
)2IYHH]#XBGV[bMKLI>&2N<(88A-_RZN^^E9?a=D9^aV^35P#AaGA36WL&]DR8-+
4KfM]^:))]4A<IR(O/YKZ42#9O(MV\R8T9Ib/GQ1.8DPKggVIQE1.J;H6.YK+<)E
:b3_G(5#58U93)&?g=Q^ZC@B__W_dK2\TXZL;KX?T:OUU;Z@FT[=:>V<cLB\D1_G
EK-LVJfIK6Nb5K&HV2_/g]eY\7F^Q4Z.<e0::^:[f.bF3GVGR1W@[_Ug9ab;&\SI
HH-(<AfKY8UZ[8A/+g249@,ecVJT?3,]?FdKKF7P^Y1[gX(cLV:F\1a;_Cc2Md&E
;6:UL8<JBNOeO\CL42PK4Z/W6P&dNa_B,M:42g4LgP0GK>M?:b7d]@_S2X[aKeLX
^A22U1<S\,g5+5<K[,(2Le/.8#?5QX?8:.Ea_+NVZSDQ(4C#ETe)+8gd=STPG3[C
S\+)T(682eH)BZJ>Y0_OE:_7]e@/LU[6^97/\a=0c&MSb9(;/#b<@M2=L6[^@HRO
&e)D(S:e]EAb&Q5\]S&1JI(44)S--bc4ASJ?+H@:GK@Z.1(dG&a+T7ID4a(4b7DA
NG;?4>3+8+\;L2PE]/3>fc-)S:f<(Z9E^9-@N2@-DZL,;^G6&+^OJ/^;.-@P_J_e
K<Y\)eeES-@C76TUf,P1++Zd4acNU)PY7=(,1#X[eC@:1e(0]^G)AP>YCf]M>=3;
1-<M>GP]K0RM4LBL_]-WHLCT>&W_4BW0E-WeY)_C:6O52/8P^UMW4NQ_3GLg)a,+
+U=WO0?,H?G3W4<NdPBC(@S+2)ZF>-^I<8efF,8&([(eA]:(+gU^(gD6>EU+Pe/#
@1c9=VV+D0&KQU<0L@OCaAD_&a3IYN9?9]?dT-dZ^HaB,^4W0.FE=.DNcBJ;[7[=
3?<abIV#9cN;D=[:KX8cg#XTO5Ub/RMY+<<MY#3F8AZ]a8/BQb=feGb-a6FU=\V,
MDG7/36=2S#N1S6_gC;Vg0U.7EXP?@08WN<bP8WLY2VN5W&2_1IV\2?S&7[-\8;H
7He6RA&3VRE31XT[68QcdMP)6I(S5VC=#IF^@<3X)Pb+ZP?@YKH=EYW,3PX92CgW
a2[.<QHRD\LH:^&E5Of;0^,6UWOe132#=MPV5Y[>+S#O7U2CW;.DC^89>KJB-=dH
EF+4[_D7IY<27XE@]Re(VTF/>30Wd/58(M>3]]CV+XD(H(TDBQa4DOdPIG,:)Y,8
(E)4K3F>US&P\8PIXLU2LC2[aBK[60;;2\>TJR_B1@GbX9Ue,@1#OJKN2-<FM#N+
GSAQOXg>?3d#+F^K.CZYF:2&ab#.WdKR,aH#62&aO+L>>.eWJ;N\-N539#B>P.X^
BN+J?,d0[#>Q\E=GUI\d,V7EZ,4^b?.E29/\N]MUJQ6^MR(0M@J7N6I0XR1+/-]&
>86R9_20NG\UHSCa7Rc23#1fA:f,I.:OW+NSO<1X]?#^7\FbP4Z5Qb7RUDc.C65f
JZC?7C^g[G_I60#/YOK\OG@#1DU#N>WEL2;>BAg=e+R]W1T0+,]ReG:f\[^Q(8;,
@H7WF>Y+F>Y_=/bFG@XO2,<3d&67>gc],AM7,Oa/9^^DH(GT4)(JJ=,5W5+)ENS2
?<10I9368,9:15?JB_(-)5eTaMM0VM0^(,f(KZTV#@.W@D#L4V;@<NM0:T@Tb#IA
:baV+L38B9#LWc;E;D@8QD[-O(2KP:A=2SOYKW,ON^HEE4Y+@I)+M])A[gMC;)HC
J^a_J_8Og/8QNQ82Aea82R9;1W?8EOdAJ4.d?F:J#)OH7d_^;&1c^:SZQ7&Scb@:
WLWY3/b.,#c=Q36+X.52B&R;M,cdLEP[4-8R5->[V1FG)20&R2>>K^(#/^GMM_4K
8@T2S4g;3g]IB6c5M_:S_(@)GW:75X=52;1aQU][FG.d4U-5f;0PbHT>b2<Eg1V#
BN8)M&97-AP;_c#(,SbC>a/-04a[aXN?_3-Z,L,^W8@&98T3^<e:^3&YAXY_7:g1
[[XebW>+TYP2d>_QZfAFW,4F@.>ZMgOFeAB+@+]I4R9J&98X:F(LTW8WcCgGEBTK
NXP+69ZXLC?H#-OK?L;2A3,A\&5H:ebG0dC,72\Age9D3FK&Q4g;JNO[=bK8Dg4A
@4BWec#I?10d<?e9(R>>J5XJ]L_C,+U/FUVV0;.^@_,fUA>>GGVFg?<_;>59W-d&
E(X)IaWB.^.g_4.#?.0QMVU)K@&0d?9g;WXR;,9b/e.Eg;87c#AcLEF0;]-1G:?A
^>&X7X:?H,?6#2+CYG#UD[-73Qd)<CA7e.a/CaK-A(E=N5=FDH)9RSC\8EaP<TF9
(5dAEK\7[3?cK@U6H8a=3O_1?WL(ea@X<]5VG,;fPS89U8?2c[=4QUFE5aH67BB^
X:S+\N5a3\K?KSDTH[A\D(NS=?a<-@8Y>69K^>VSB<E0OJ7U&&(/J^Z[F2^eace9
MZ+GBUf3.?Q7S_+R(:&Y.K<&f&(Gb):\df[#-dcdF:b7Z[RZG]C/^U)^@@)2L@fO
#&TTK/<U0B]B-VL;4:Id55?-4O+]GFS-DffWT],NUfVJL4&/F&X),X#]/HMT(33.
[S63T_E0HTdK518b9D8(fRK\P5NVRE5:=TAg0.?K:ZBaAPBRJ\_@eW_bX>#T>HE1
:.ScW3M1LId:gHFF7X42A4b4:B/1W0-M-+fQgS<5f8XT9^;7Zc_<;/@3\#^CR+2E
PNDB\RHA>J4dA#8g8g\(a;Ga[:@bNQJ4NS)D.JL5aGR4OAC>ffb:]=7^;]c4,5=f
TdX.=AR<Y=]).Q_J+1KbebG)Mg8gJc5R2eBHa[^_c\>YU/Y92:A4RWd\585abAdH
B^3;/IM[+0#WW[T)\?W?K8XTcFIdUU937gB[6,&)gV2\EIM^G-3\OPD:XdU\=g(-
7;Z-H0HY#@=DP9219IN&-&4dW7>S)Xa,&SX&;^(39ZXKUI3?bN&-V+5[^2;6J6LR
>bX?CV-EG1T;fEK6)6L.9.])cWR^+d:.PEg[88:;8f\_+C-2XcENX3BYB1?R(@-;
JCCeMb?4C=3MA6>NQ[;32:(2AgDY&89]L:@^(b>^Ga\B92N-c#X-4BFZf26Q,WM.
H&QC.T\R09]<+Y6FW<>^3J.GJBVb)L>99EcK9AL/_P8W8M0T&W5AVfB>+_YIYI:B
T./+dc.eSOCIX0#[2EQN]b7B-J<.;Y&LdQ>#0MMbB::=-#VEU,;2^RDTKESN6_I,
g.EBefTT7(I.^ZI0[0#KW1HVdC?@aaEP1-O0T3D07\-[I3TLR[R2:(G65-[<;ZG^
?d3YRR;^1J#CEIN(F_^?5+O2;SG8@5?HWM/_29+gB8)b8-AbR6QIBa(#]3I&O515
IVL_)&]OcHYB.[M6=1N#MP2f5AS6&1BME=c5LJ;a7bS(4ZHP-7EaO#?_2&C3DL-/
T)9CEZ=]NNX>>e&@GN8<3,#+S.ASUbSf_J^5)IN)H&^A?L_a5Rc2MB8GK?S)#OR6
)NZBULfI9<RA@_A)G_6DBIc<0EgNdSbI1CQ&Xe0HZ9(\aYg4(7([dNC&)GfQ2>I,
=(V+\?IUgH]>dT:2Y@]W95+SRe)MV9dSbSWVV)6GcROa&;RG-W#>1Fe1H<B#eE>0
A.4&M6LH;\>H;WdS/#^a<27IFB+J1KP[a?5(bO7G[bSY2A-0g2[W[Z]+\P8>>MCg
/JM]BdDgI0)5);[IdXM;J?&GESQbF7HA4WU>F5K9)RcKFL)[NAe<cN:&dN8(-YS&
H&G:_ZU>A@@GLJO?gc3>.E.WFY\JF&=;^WL[cg0#XfHW;V2dM1dU;bEP^O18C[Lf
D&aRT#?9M&MHe.43#YHIQHW[S#@dEX6R__2W^8OD5+>GMfY?d:f#g&ZdS\1cR^@>
9I4c?@Ob:;&2?+Q(QENXGAD2JK&-?F6=7IOEF0W8A=W.P[R0-V7K>f@^+1FQ,,[?
[4Rc,M<>69+f-I4gH6U>^E(U@bT1YI:N^OR4JCcMMD_&TfN:VR2Y(88+AdQ(,-S\
0eZ4feJ4>H([b?D[]MMX0Z\HfeTY]#U5&/PcVU[OS2;(=A+PCYG]AK;9Ta-S+dM[
/:\g4MbeT+H\>MC1(29GDAYd)-I=dMW6><=590?PNG09S/KSXcOI,UY18bcW0NgB
\03R@Q>&aTcf)bUVbYW_Zb]L\(]XT(RZbdXUC,,L_@H-SG]1dR@U:9:+4Ge0TS/1
,\3ARNe2FBe2J[M:?TfL]\8g49Udc1TI(VIF..Kb1QP[]YfRH&>4VaCV&6+]KaHQ
WBLeV.8H+8H[)1XgXX[D\JDPU^)K=&2A4)3Cb&+H&8NF,N3+f[g-_\/+>2fRa3OP
X[;F.#<5L(ccabcR=XEWc>,S)CAe>1WDa12c5Y9I)Y+F.(X69NLJR2H32>9<DX@I
LI[-?;SHG.T.=ag24,SQNWG;faIP_^7.H.eARP5WCJDIS4#74HP<ZY\EKR2fMEW,
UR[@LfQ5<Ua)1V@\61,F;f84+&.QY3/YS,/.:eJ6A\SW)[Z;VA@V]T(/Gc^R(KA4
a(c^;1&8:g,IU9G5_X?AFROaZ;X1=)9>U;>>H-=d9TZ,\^BMd;AXdXU+CIa.PAcb
cN>U4c6;eVT<\19224)#](?2_Z(g438I0]NN3#3Z:&dI3A_^B^W5_Pa:e,DM(?I:
;gPW\)R@U,c@Qc2E;UfKB-FDUE31^=90G/WF#.]Hf]OL8PPG\SS.;5-9[&W3c7V:
X5TL1_eG^_EV+-EFE102,CI)93dSDVeYP4G0Q^.OUUc=a^QXZ9EGIZ6J-b.HOK0A
XTHcM#&:T_Ia:DK;TW>@2EE[N51WZ5:3XUb3bD)P7J8UQ2M>ff\CX;Q#_C-cG5de
b16&7_f;?MS>0=)E\3CbVb<5KGC1M\+1f8>JW-2^H&WH<_[S/D^LO\&g:9J)1UD,
3[?-6?Y45M^?CQ0gaY,AD>3d@J=(OgQ0d_>6MVH55?a2QN/1aZEY[&62F?##SXL&
WfU-N7EEK97eMMcIW1LCY?KSTY/+2Z;VU3e7.Od&d8=8g@#L0LQ6]5BFaYT/7=)P
3A5\]12@1H)#&f[=M>cKdB\E)T;&+?1[&XY#J0>(E@)c39LK(XB-<+4PJBXUd>O4
a\=NOH7^Mg@(8<UKBQ.MVY@OCR]IR2ZRNe^3d:Hf^bQ>XI=^B<1dUSS#c>Sf^e16
JV3gQ8/B#,]U6M<?VgN8>LEGaZTd7b7DDe10E>\8ZB50+C>#g3XZ/@Ab\_88;3;0
R,E)72D222[JHVdG8.d#VQ9f>9A(=R#G&Y8FJ/L055.=@/C27]b)FT@FZ9\(d@=L
UfVY<6KL+]=^D5L6Sa76=IXdR7Bf.+6b+7+HZ^McUPRW^KZA7.68G^FV[69O<Df7
KHR_CX5UXfBD]17&/_:9[6cQ_>f]_KaYY,B748X^YSVUJMZJ)@M\F(g.eG5e\_X0
1?UdK6b&>YWY1?HcUE.&CdY4C(9KbKGB8-B+B]Ae[ZZ^#P66Z^1@>9UeOEN#4e:]
c9Jd#\1Y/YR/8(/.#5T#WN9LD[aRSA&DM)(WFQ_[IKdeTLDH^V<.a-fT1(+O-FA1
<@H)bPWF,&13>WRe&LI1(&R<,7KM[[@_#]N9EJdD8MReG]KM(Q/WB61L-#][7Q5T
H;YXd+?bB7Q3<&-DWTb?U?e1\Eb.O:758E79+T/e3CNJ0f_,3WPXE>WR1,L]?PYW
7(@3W@@UQNSM^&1/L7,Fb8-1cg2W.IT7\[?P#.:\/A.6GG(]NYYE@Y<Ug\[e2401
fGT>NU7gM0-DGW#P+U,52QF?X,2,c0V>IVB_ZNfO33/VRV:WFFb<]47)_>_;]d+;
dAeb9KB/16D3EYgBaeMX[)[a/3\^Q/7/Q]R)BQIXcZB>AWcA6M,-WBdI@3=TTJ7H
B=ELM6fCPf,a3OaZZS_b_D]gD3_d/;-\dNR8I09NPYGbbHDFN(;9?L?7dHM),W&F
<DZ-JH7d.UY6GGUJOK\DK,<)1a^##;6X4,2)T4BU.8\Z,G9R]@/ST\B2HVD-:,R&
Ld3@,&](7BDZaG#S1b02<RR<D^A[Wg5B)QM[_bUVLTfgd-LeNW]gSC;L(+&]+D[T
b0[MCeQSR0;MXQLV>J_135A+)T\BN;-TK3f^?<_@M#389&O38GIPG3WG1OO<D4(K
)K<E:K;8RgRQXBZ:YNMeYeBQ_Tcb#Y_&3D,]L&=gIdbWB<+)?;BcPJ,8f\HYO5f6
E(O/CdPT>bc>PO:,?D-R@#K/.L3+3TXG]Z7c_#9&<E<>Z[V;f^bX7],d4g21<cf&
-O<H#[)FWaN9&(76APV.a2?X+g)f5b2(2TI,-=9<PgVF:PfAa1Y=9e4:VA1J)3<S
_Q-[c-[#.=<_PIC#XMA^4Q]=A/A^f7&f.CQa0.SP#P<^XR][]CdHGXH2H^\gK@<D
^.3X(?,6[7cKN_O:QU&0@,>V9S5gE9^WD5P9\<W:]1,AR9bAI9EYMQ+,>QUFOZ9)
^/;956-32\;b0=\a]Z7HKgf=^##R0W\8Fad+\LL7+(UQ)2Rg^I]84<.XV2##.-JV
dcKZHg&@HMN(=7VAA_XS-F>:)WCK&HRa;B,&dTQ(E/UW>5YQT<YbO:1E/89NQ23Z
^;I8)JE#CcS1df.U#eDE.SbfAe<D4O,>?M@8G7<8Z8@1,/EeNP.cZMY8+J_]^V+#
HeJ837B/:8<+6LSJX=[PO&GXQWbE.<T]Y#)/^dB0YJ=L3>V0&_1c&0KTEVNV/>=D
DAZ-[ff/Qf+A3bg.a1fTB4(#WER]4Sb644;1ED:EaeA0X3J4fL<N_NW<_FaO]7aW
R5g.W.]=DO)>-D:8=)GR]H8_c<SX5<U:X@_;UJ#NC2+)7Zd]aIP>?7D-f]gZEY9X
<UG_^ef/]V1F9=W0:6ACCYJ4P<:NbD4]:Oa7?5G&#F;A56JH,)e47G6Ef]75/?g.
&&.X<P0QSO#SG)dEb_Z<>Z4BA;<6KPZ#ab..-Q,Y1>BAA+_5^WW6;9;IVGEE\FK<
FNUX/&YfQ7T/LOa?9Df+U5G.A,NA.8QXgDCC_H9]Y[@9/3YT=e[M9].9)c?\Bc(;
=f?NQ7Q5&g-_\\M-O0d^5?L2Ve)>Q(Q:?f46?#a#J-?CC>]K3AG_2?5VA.T1#E\6
X(&g&EE:QG^;P<X,)eA_51CV_YSD.5N.GEQB#A.=?;4XJb+SOEQ53a5SM/FC;XJO
Z+c.32(F3a2SCLQ/F,TJ[)bHP_]IKJ[aS2;9HVg>/JN]SW\V6+N2;8bc.9N/9=dN
#S&<1T=VM.,PIAE,FGQfYP7?\L1RTCWa>ZgXffZOMJ,Lg#@AcB)O-+TYTLR2,#V1
SC=\,9M01UAg&.GPA42F=HFDADG:3=)OG+EbA]egP_[-bPFLXd&bU<O9KX)F^ZB^
^b?8>&)IG9.-5MR@Q[W9=T08;CC#PSYg9YNAE/eG^WfUQ<gc\G:X]LL;TPIKT^J:
Wcc_]^26<8TP0g@e&U;8,VQT22CJgKSI&YA:?4M(-_cT\>L/fW]/JQZJ255g/AB:
\^P4RO1(7fR#^Jf-7M;/Z0]5_RGS[]<@4cC4fHCO8;ZPWRS;UL_UW-&8>KaI7\:3
@3HNCZf9eH43;KB[V\B-]KDdZE3DA6g^Me]XP<FeBe38[bd_JBg\ZG4Z@PFKP=T_
39K1UY#0<YE2@,dE:[#/8D]Y+S8Y[_,B@b>1IH<:60^[3XD7/39\WY^VVS+FR#0;
/Ja-aN\7]g0(ZRFaQ#CbHK0<Ue6S4_R#S^Y]E]aBALMFeUDeTVd(<&P<Q>JJUYW)
VURM5Z/bdg\D\?S4L:a_RcC3=,?ZO&H0C(;OS3;.c)e>2-##8UcPUaCS1<G.K6AY
A6\SW[N.[GeC=[KFJBF(EU9b2PO8beS[O0GH;UQAMeV:=,)]@8W&)g&QBM]C4P+V
)NV)S\Sg^_UI83,\U@(Rec=FHN?6OJ?BAfJIe/=4Y<H0_]S3/HXI56_CJCbL,1WE
P34WWM4Pg^2Q(0LT4De1O\@<ARD>Le\HI4eD;LK[c/6f,J8FJ0Y0+\N0Vg6CX&)Y
Q<<3F--OL,:INF3J=K]8QHE3_N=.fMb?6JXM><_=]DM=<RH1gC)VS]e->R43H-+R
@3?4,-VD+P<eL-_XA2=/K(#cL6BM;:;P&XLPM1//X?A1McO->K8,6>EJ6F-OUE#)
e6&6g]7MEWLdI-/IS\Z19#.2;8A59-A1:5/UI\c(eY[Z,WGTb2M\K07YE(-eX2P9
+4fZU68bWRH7CY8a+e8#<6(,T8&N#&]\1fF[9<9,9=;8-]/-O,fg1.SR8&ES^MV,
D[/,Rb-^9S6e],RG3]S335&B:7>+-24OY#@-09CVISe2,P(I5.)G0^JOO..L:D2B
O.-Td@\9D_NSOLM@COWYRfVTac(_[.9=9QfTUGMeR+]8c[_@ca5&UN/YA<g-g0d:
=G0HE#5][69G\K.BQ\ecV+DD\AH,)YB.#->NUUS^MD2=RQ;0K0LB)IQT__V>90VC
@;W9C2f[I1H+[.O?ae1-dZ9fe,UE]CFEdeRTFb3dE1b0LX@SdPXQXBg<L[@20Xb?
9a1D-L+3@Z^V:X0.g1gP^?D>@1NEYJ2RH@)5Z]9YU3::BA?Of<=:^XIcOG19&@If
@A:MF/e&-]@<(/QA1DA6U(d0Zf<4B#@C/-06)Ia[fGDQ4.:X9WfTbW\SD4TY^<CD
Y2=)KJX1@c:5;H8-_77Q@a.]175dP6_fGC.GT2X;G/1+R&e4UA[A1@81YF//^./T
5/9Df>;_>0KKDKT5@dJ#9.ILQLd#]8^MdKE=;C:,RJD^a^>O2d?-23&1^bE^YO3b
g)XbZ7&N#1dB=G61UW7[V6(9G9Ce9Q?K.>eIB0CYA24F.J#7GV>@db9[\DMH]#MQ
NO,?dG..-Z#O6gf+eC+P/L?->;T;@feKB;LB1)bLO5M&H7+V<I6[)I4H+B-?.Qg_
PMaf\cgb&SeNDH9ZgGZ6(YLCc7DDK0HXa^+AN0NM0=VX<A,X8U^gYUC8B(XSVS:9
c8M5KdgLZ]d>CG2;C2FQ9GU&[H[TWKFc>HXKWP?L2_g=S[MKG#g9KgI_>\/d;2Ze
.FCG,<@ZU?RUTAJ]01@WR+>\eg3A#cA7U8FAIO<3?U.EAT?gdJJA-/0]K99V@:1g
91d]>dfH/6:_.P4ZG\B&-]J\/^,PG9OG527N_;eH<SG2[3A:A=I<.<;F[5T3S5?K
NOLU9>eQ/4Z[0))-c^,1ZDMD_d;8SE\OagI/.,<LYNJY63LfWE5NI8?J_AEQa7e)
,00Z;._B0Ze6bL,?79+b>H3IX,;4Z,,\B9R6e9,LKfU,5g5B:NK?D?ET#7/#B9P]
[M+Q9;O_(B1RV1_:0Jf&f/(D]=I:O0dP;PBU0)YHb1LZ)JdeUK=AA.EBb#UJ8YEg
_e);Lgbc];GTabJ?G@Ge1[.7T\D^_2f[OHK#1O/?-=XR3>a5DM>B::Y^?30DC12F
fF?P/BQ.:-V<(g@VdMI#9L<g+A+18F.L/.?fJ0=Z2gE4REM]:](=;G?9_I8EKR60
2c/MQ&A@c,N3]?Kg4,=;^^A9BWAB9961Oc4+>6(^8/>]FHeYe0C6e=cEL()^Q-^W
;T_G)I)(7_1,H]@c&eU#.cPCb-0dZB+5gG2@DQ9&FJ1].5V>Q:^;-6UK+J2CPWP9
/@RUV7cDSU0EE(geGFgU,L_):Z.B7M(c&g9W5/AIIe/APIf>MEZ2B9cE>E^8)+6Z
/ZT3^ZD.#F:(_&RI.42e,8XGCcCCEGRf\H8^25Q/\Da#V6U4/(H.1?7.V63G^W@E
gCCMf,U#/61[Q#;&85<25b3?B&//4IdF]d;_:#+8+T8XGA.2&V=<IN^_<e=EeR<N
MbF4<&1=MA&@LcJg.SVQR/>ZJ5f3N\:_,9>[6Vd.BH)@[9RHY&dKYb8fZ9RF0D^Q
1,MFZc\(:2IZI/L)P;1&K9AU6]f2,Ag#&c-cQXSY/6c#\8ZQeP\eQ].>WS[)4daa
g9XEWaDH,06Be:,gT5(V2+&:0B4bN>,;]Z+T:_\OX2J58.g+0MfY.AIbLN3V\bGJ
B0KVXPRfP=?+.N42L,c2^2//M:8C6IU&9?ZfE_75)<YNC52f]NVcT=H].EIe2QAB
HeM2=EJQFg(R;VK[SZ9<TC.C((CLPOf(bA(I[G3LRW)QVYM5((0K-8ZY[N-Q7@RG
(9TA46=4/JWDNDOURN3+.0M3bEM=HdA3:f/)K3^Y]T5ZfSB4aOP=ZA7gRAdS3O0,
)7KQ>__//#\+[BCB][]OG;PWLfIB-b6Ia_SOEN-K]5#RfQU[?/AK3;X6H3:0Kf/R
2#CTDSKaX&b7cJXH<bC/U7Tc8FV4SGV^ZKUIM1K-@IB.4@3(:CIg[W9:[T^(F4VG
VQ?M[;A;3g83b;K^HN\-A<e1A>X4Q)c]_GUN&)/YEY6APD^bgS)?;df15^,BbJ\5
[L5gU8QA871HGJGCR_^&Y_4AHb#-Q<g2G#IU0MZZ-\g1PZe7?<=+@Y)9;.B&.8^=
.P_B\>?&aB7MQ:TVH[718=35dNA^Kb:UJBRDbJgMYFJRaC2]:c4D/J?NZbUQCWBR
+^E)bBOHI:B<>?Sdc1V7RFe]-Q;2>U=9=4cSK4B_/?BMXT1b>@K#_D]]QFZNc_,M
Q/63].AC1T)7/??-(/3;f=QZ(<QZC5L.@9JgY-.,G\@?feWLeG(7=3W#P?Jf;e+,
BUOg4gW&aU.K[Y]<Rd1@,a[9+dCFTBL=ga1S3L<K<f[S=/RBZR/a&IFK=0_[X-;Y
TEUG(2b8T5[LOT#]e\VS#(B=1gfQ<PUeReKdZgR3G:7&Eg4LJR>[G+#[a)9Dg;1S
R0-XO<W\e;^<F[NbK,-PJ=EBS/0d.<G1/VJdc4(D=ffeVEO??e79\J/S+:&CGg??
XIc]&2af-1,Y56ePW[]B)=Q3,A.@.Y)Lbdfg=76ME>^aEJ-HOA?9CGg=BZ7+Z#P^
;@XK499b#)BES<ZCOKY_BJbEcc.?@?YI<6Jd\O;4W7.Na_7a^bL1Kf=.W?4INQ-V
O<=.XIX(9/.e=;?Oc6<-3+/JEeD?ZF[a/=,>,D33XXG<eK)a/S)+2<2,#BR7TH@S
NJUU(@9MO<HO^,C=SC???SPZ<;XK(VF76^M/3TOW9f[]#?#((_OG_HWI.(E[_,5\
U+eIg_9+@=9\6I)71f.V;;B7fc?#,^.B;XBgXL:b:UYQ9O.]-3?IFX=FQ(.EeG.8
7)_.IA54O7R,0R-/8NcBa>@gMDgQX:fVJ#C52(_a5:T^R)1[ZT_IK]D^83FU0TX^
R?8W>bcDQSV@\N418Ka:#(6K23JJT]2d<FD;:PYYUD2>Hb65;_-_Qfcb4)YPS05[
U/4=e>W^Qg19SHG_e/g=,++L#.Z?8&fdO+,Ce2E0MR6#,Ib3)DN1@[7/_Jf+WH8@
-@EQ5cP5.6^Bd473C/gYOC0MK<D<ZC+dG=?75WWXEC+Z/0BaZ:S&K4gPIQ]^DcE1
=MYZ,VdF&<QD__AOW<YO+(<[0,3G^PD:fSYE,DVe)d+00@854XZG5B69^25cd.Ab
9aR25Q,NQ,Z\EKCPSE\=JVc)-Q^<+2(IaY+2dBO7e.H?98,4I4#U&-,2/d(U_/,B
aSga.8KdOHQgV9X/>X<Ge1,0+8U\T.^H+LeNf\]A4=B/@SV3eW5;(INZ[_G?+#^M
U)NOC5.F\W#\ICH^W/<#+)?+S>VHVc[@OV2(/DNA#^g.75]_&8X5IB3?<UBD-2<,
F-bR^5ZQd(91\ZNBX6>e&40?]9E(ESfHMQ)YZ,,^3I9GM,FLH(#-<_@X88d]+bR\
6Vf]9YT?de.S006[]]9L.O3U598LC^#)+PD+3GGM]cc)(R/P81c9Pd=@^/VF<g#V
C<cX@/?QVbTM6GL)Y2a#FVEbPZ=_2?2F9Lc8TJGVUOGP\/4eK80X=):e;M<YZF35
K>,SQDKIQbdaQBT+7GV+]TI\NeWFG0b2KY0O<-HK/-,FJ85A&=BZ[=CMWaZ^G\,K
-^.D#97B@GKLAD#c_-1+SN.B)ZX0TCAfIY5PIW,J?7NBJ.[T(4^HYUZ@O1V@B\3a
U^c<J.a6gX[+1dB)Yd:5(XA4#A_B)0#HO74,gL=:R4[+MR8GVP-fa&3YS>?S.Gg1
Q5e),ITZ:c2Z/EXAQNS=T-P#<-@(6b</>\Y.B&3e049:,@<>[d\\\HIEJ&;);YY[
Z[3eWSY#d)H^;Vd@\&+;^a[AGSVQLX[K^\2Q3>cFVd5=V=QCHQPS_:3D49<5MJ1)
+Y:-fS)<B[gTg4,M+NdYG1.Rcf6_cA39X)A;S#Y2?V?HQMW@Y:\#M?Q[g68SF0UU
7O/[Dc4WK2fG&X+/60aVMgFN5Y6VVDU;0[AJ]3_-,XB]Y165b?=_Y4f)#G=KCQ7O
#2FI7Sf;D7,HXVEZ25T@MJd5:<^WTN1+W&?(e,^\VN=:W#T4]+()<Og6A<KbJTL/
=FBB?ge/)3&PCK75Ef&>)STO:RQ0cI1c?FI4bNc>J1@VN6V#RE5W>A\^cb#J4&O9
D::3;-2)eIb(S5GA(T:/gU6/gU_A<._g-9,e<W-I1a+OZE2H\42#DJ6ZCbb,3@V.
f\V;#M0G5M(I[-1E^)L-g[N9-_&3B@-2EM,XN)&,e4^cd]F;e_I<LRNPg@DPg(C.
=I]+D:1G=cFd:J-^dZef<4NCQZ\CJ?5536g+YVNE-Q?]U3g,C\&H/dV@QT1R7]dD
#?G/aX,JC\&I[SEY?Za06;(,dI/KO^FRS93-KIRfO@-@c;S4EZ7E=;&(@T2IG&^b
d82L[6bV;U/7K?-E<UW^QW(Q),.fOKBT?gS_e&^P57Z/4Qe941fHdCO)J,fS3Ub?
4.VN]Q#EcTB304<^0J[fB((F]VOJf9@H(DEf(;POPD+Vc-Z/3H584<M0-NX6JY+;
f^W7+2I.&50^cd?]OQL23#Y^E776A+_\NA3(36,eXRMd2XJ(DgSEIK4P2b=+=bA#
XbJ(-,VCM:/a^.0Q9a(6]0L>B&Y:I4(-@JQ<a@6gg#B]_43.C+.IF680.CGOfc=d
O82P:/1L[?.<^9]-XMM(6?LdCPb;Y,,:F+7?&Sc:g..(Z9KNHP\9e&&=O59U#G[3
a&\M>\(5Zcd3PZMMSD;W8&MME&\@QZfX67/(JE+^gFG_H;V15N/]L(D#.1gASg3&
\cI]8S/>e,bgA+]f?b.daHBWG<.PJDMB>d8.gdd#&1GZX+HFYg+S&6PN+1BRRS#>
V?1.N7A+:/H07+e<887I.:]_NJAZDf6-8I12Q-0V.cNZN/>LA^>A3eB2-YId/DZ+
1[T1ObB^9Gbc;\A.[#7J??a(]L5\ETAbe<)c^OgaLV55-9f\J(M1@GLA<VeWa1)I
fHPBf;1)K@dYc5g,FY)2UM<[A+6F+=V&\CfJ^N+Z8C6Q)_GI?eD8,>44B4Y)g)],
):I/:KVO^L0]UY9PQANEO(6f+4:1?Z+0RJ77RW65#T3@b>:TfK&a3d2I+Y.@7<ZQ
.=f>2E+2.gRBZOJAXMBBBVR>CCZb^+DWPGC9S_I2N,:N.K[/R<W9-<>1REDb[(f;
ZGVSUO9Y15=+ENcN,0G?UOL0Ibd^SeT?T;)a=L0=df>7EQ3+Mg^S[+PfV3R72XM;
UD6@YSbEX@fS^I?O?bG2#WTgW:Q<5DC&_V)?=&\1?V&B/=77M5MVCYG_\21^TK6^
TM&S#P)EZ,,(_RbEC2:3C+.IBgS]2.I,<ZA/fGe;R3P(3/]_BO5PY,<#<;&/6(W.
FEf-:BN4=N&,@1Dg?X4DaS:_Oc4+M90g6f@&G.&E9F0--Q.Oc2#85T)0D9,,IgbY
a/PDU>S(V7#=,[S<H1HfbU][TE[RR1AE7:;S50]\GM=2+)_eU;\e5Y5_^d@OLgf;
H27?F4=RAc[MJR;>#DQF9EFa.0-52cYV-a-6+S__Hd:FL?5(#M(5.B<DCLX15aCB
a@V2a2==Y[=?1X#_-ANWWQaa-f87K++Id09^P,[dW;Q,91G]/+40V/=7]g,Lc;YJ
+MF[&gZf:NI[65dK:8I#a+90[JIXP09c;E4E4QMSdDML8:;5V,d.&Y21-6L+6Uac
fHaM?D33U;\O9BBCf#4bP9M10N_,<]d]N2VUH?7=&E)(A7^0]b&)FB#PKL>MMf.c
0T5=FC_Ea:gU74JYZ;aLf9=,#NYOaMf]OfW2U8FRZ4&(2RdZ&Ca#@.V9cHJb@cN3
FRXI<Q#V=37)EZ>8NH@,[)FC=EBM[G6.Z)=Vb[b]R,D-,FXTaX&OC-1S/#_F<4-d
b]3;V75S)TE1X;O8AZSW_+/F<G8/0(52@9/OW66T4P_E[CdWYP=)V4W=&<g1DS\;
P/bBGI,?)-0c>]K;b:=D40QCbY[HKgK&-(>81S@fSU1b5))(8NRZZ]XUKIF5/0-&
4Vf&UCIE(WD>7KYTCfaV#W?dHF3NDNZWY\(+>3_HDF7=Lg+_RD29b)J5fMdK42L@
Q_G_bNH3::>2a<1=;I@Z?6Na3#+DM5GABBU/bN#3;J72@C2FOQBN4VVD773@6a#G
]>d;YK[g:#XO?WI/X+92D@g^MNDWCS]H0M_H/<Y8ffU]Jg5D,TFS\.BY^Y4613^E
g(FCPS(ANg(G.bUQRXf4.N9,gfT6P.b3K787Ne@=@C+Rc@4^6Kb5RX[8:<?WC@,L
[I_[BZYe&F=I;O25FJ>-_?QQe)W5N\=K4PXf:7gfS\)A4>AT2aEca+c0<1SGVc6(
Z^dc,U;(BY-Pe>_cbWGcb5:g1??4<^cXSf7B(2NZ<f<2NECJS#.7^[\4#-]B,GSe
TNf\a5ZSMe-4]+cI)_B#;6[JgN^>N-8V8D3G6S3FGK9YS;YEReESIEC@1E4\=TRB
(:)C<#Y4ZX=A=bF]9R7(XDE4P8S2eL+UI989N0SLH.<FcP[CA9Dc56GS@@U-F8U+
/49a=@C,R,U/Z@5_OH2fBQNDY\(+XU43)^4<U;96gaAUQ>Z12GUcace3dY#TOD^c
[>RVA+_()VWGJa_KO\)AJ6-DP-7U)TYZH)SfVJcY&Z<F;:3aQ_b;10W07Z@WHgQ[
SUg75&cX<=8K[Zb;340dDLdd:2:>d5AMPL@(ZJF?,KFN5M2<eLG@bgF1R\H@JMZ9
Q\=9FRQM??WW?bf3A?ZPB8U1aSJXB^bKXQMXB@6]ISE+<LB<0?&>R_SHSO]5XTLZ
OZ^FW#<4GfYZg1&Icd9>>([BeY.^Y^E5-?N+c(QO#UbAUW;UZB,R;73a,,HA<QNa
5cTB^1:)Vg<)SRVEa&E\\R[Xb[UY&=G]\]@7QK-_VIHaO+)O[8Y_EeV<#&I(XdXG
GKbTT8^<1DR7EeR<,f/,;N:R(Bdf/0B4#fJ8:]]PQ>.;/&OY+CW.CH9ZP6_5[DeK
UL+Zb>;NPQNgaOUIa^Va+X<eD6V8IcY[TE8>J?[21SZ1=4:M(EAWG[2>MRZ<I1&)
LNR,g;8W(6MaL(fSgZF:Z0LPT1c@f0^P]V\R+M\a.XeT_TKE(T&0UR\7CMe<NYX_
VZS+PHXdfaK()XeXV;9]T,>QEc5YJQ#PNLV8^<1L4EXKaYWQ73QVFeZ1aVI3S/d^
4gH,:R&458?CZ(.WfMSB>#N^Z<;dZ,2[#:_=SG<VD\0RF?<-/TK,-K@=#+Na0WK6
dT8E9@B:M\Ea(CO@_eW5?06XOPDXIP+R[a:XL7L=M0S#AIcV:d^P50?2K(a8&D+5
QTV1W6-Rfb:g_>)#[S<]b)K3Y8V:gb?456=Vg:D/4^2WSK,6f(8S[6:0[=37YG/f
5,+_[3S=G=G8GH=VFXa>QOEI4_NBf^&MVJF7a5KYNVS@a&;#_2HGg=g^2A.G&4&g
L8@.d?;S)E<f7132H_CJ;RU)-FYZ<M-&#XPcLK5:.,<O;QV&NF@0IS.Id/FRGaG5
#:032-KDC0.cW.9D8H:O@:D>7af>9@Q0QK[)#Da><Y.NdI2,aa,DP/SU#=WW69#K
5F<T1H.-g+G&1]A#f1@<(IA?R0+ecVeVS+eL:Y5G\g3<W[@M(P2JE7:]Na-d=VUF
S1)b8<e+g9Z14J)E3;)=Q36Z@d3SW&:AKK(e5J+7EZA?OXP2=27cDR&K:IR_-_;4
De90\I[fgEbA-CQbAOBOV9B?J_1;ALA\>MVNXCWP=I&fcZD^,RI9:B]-;,Ce/4RQ
-BC712C],8Wb4)?_.^QBNE9L6Xf(DBX1]<)RAM?4bb+]1g&\5\/>]Dg&bP47fRc^
OYA)4M8?OH3[C9_RV(3cYL13VPB=3)T?V^>/[TBe[/R7<S+]W[6Q4.CJ+c:8RL48
\U0VK7V[@\U#=FNeX;N#&e6b51a__H-CM9SHdNe:R.X&><ZK)Y-G9L4dS,8G95/G
N,PTSM@A?3gV4@c+40[(UU4?2@Mc_?MaK9SSZ1?<]_:4SecW_B-^;]E=GLT;9Z0F
aOPeOOOOe??0DCG2N:eQ_DFG3/+>\dFZbeF#ZR2\KX&)4RZ)XW^1E.;f6MPXNT;-
U5,)F\WXBHg>fTD=:MVJ:dO[d34:N21(VF?<RDZHZ0;g->a7D80;Ue>7O6I>(6Xf
N<-U#;8697eaKMO(fbR2U2-CN-U(f>SCF]B<dBQ)(RFcS-:,F.5,>C)B(8dA\<JM
f/+NSR)ALI(W7IN/^_5f_YXg=S,0BWN^QWL^&-EDI(.cW3LX55GG-7C5H\GfD]_a
]f7e^f]NOcX<dFbLBMO@[67Y=P:[Y@LOB^Ie9ZcT]f:8Uc]b-a0C49f:gaZNR/+:
Q<)EC0GB2(WR855DUR[Xfg(B19_05U>:CYN2L(AJC)4#JMYf@]U>Y-0GWc<V)A;E
g)HAMe5)73bLWX+=bcZ1gdN/4L#V&U8U3L?\I+-T#IEV;];8-,+XOB4@_<g;;V.]
V9;VI&66RebN7Nfd&38V+,N/^ad)R&b_.DcR6b4/c_6)-+_O\eJf^g[:d?:BDL>3
MV)O@I]&_E8Q@;K.LXbLKM3EfP:6::YLNb6IIZ78.JZWF[:88,C+_DXD))+L\eOH
#9HTL?H.>.,TY-@Ec_I\44[JQUE<?Y68=XfX\T>)?X,AVgM\gJ:88\WJ@<GQ.>d:
+a)FVHN:=KRM=J[4bgd:=^/&]O0dCI=V_RMgPP=AYHZ)LNL)N<0(0W2R>M4&MV(P
>GXNQ+X\]L29]5,5)6c9&<KN_V\]=c_[Ac:\O)21XHa8LGN+?1eIa>4KfI/_L25e
=f06]c-CPLAGFA+@H/aTFE,M\&F@V=fD:255SJXg(KF;MeO4S;UNWPM@dAS^),I#
2SE5fd^I>Tc,d@=^FFMa;?/IW:G:<fI,b[O2^aJ<QYR[I?f-cc.2Y?D.YG2VFOD[
f]VOe_4/..WK?MTOH2gP@&JZB#MCYAXI/\LOKAMd4WT9b&T/Te4TMb8.M:/5K?ga
6[O4eKTY5addGg[SMg)7X3&Q.+7+(.d,CU,78<&^S;PG^eOTO7F)4b?,.+YIc,NA
XEbbR<ZSOc11e/2<JV4G?\FPg&2La]+T.X;E;AbS3Ha[8C.<M(;WVQ/(51<a1XU+
0QM0ULXYZc6MK;W]-Y8+6_<5?>ZNK77d142MDHO/HR?#8D@.]DFBaZZ_YGQd&L_0
C9=?PJE7T8;E:#eT?P64Bd.+RWaE^1Y-fI^/C8FKAR5.^&X+AW[T<-<1ELU]@]?<
FGSE5>[J,b6+(H\8]JE>#\Q=-dVH;VZ1)H8R+YNMY3DQ4(K-gIJC2S?ZIaP/b2Z]
1+>dB2=W:&^4/I&&J_99XDUECWY^>[4Nd1EOOC@9HBFB[)e)6K)U_-;SV?<L8(UF
eSL)U&2cbOP1,a]<K3]18IYeGQ#:^[6GJbX]]\46=BR1YKM+?^bAEd.L#R.,NO<L
73bZ5^?F)<L-+JeEgd<AI^#6S_]f.IT<BW[6MNLS;QEVX6\1HC@(+XS+(2U3YXBF
S>)A9XBdJ1_Ib:ZAPfW(;NgTaN_aI+<R[>&K[1G3STXXeP?f?cVL/U&g7I[b0;RN
G[I);dcA(FIZK4d&-THVb5(Jc0MX3KEV2KZ_-_]?;@R^g(&W#dY)_G--M\;d].SE
VT/N+ICHb?&@aBe5MTA.6I^DRR5>-SB.<ec[1]a(,T#\b4A&F5-IF^+)SX&&113.
3a@ALM[-9+I+@WEgT)LJ/^OL.>IDEaN-#dJ963;_SD0M7g4(]J690aWTC#6F=,e[
2(]U0AS_0]^fAP(M#2_Mfe)=GS<GDH/E_U/UVceF6J16&\;D5aPdYL6=>OJ(bBOU
P5CE@-g(:M7FHXMIV;2#Z7J]GQUI<[/]70eWXO43R9K\(^E3:06>040_]FOZGd_U
R3S/<LCa#OH<+RdeOV)CVBQNEA.8#RN9V6NO[gOZ&AN)\AHO?QCAe-ZW#Nd+]U9P
/--=g.IFQ2,D55@/ZQ)<TQ]RbMD:#LVgcJ>1X.0-M\Oc9CG1e4[>Ue3#Y4S6&GX)
6,@><@3<@YGg&F;NJc[V^Bg<1_>/:(fI,bUH[.M,.PFYEH2b1fN/f,2/KG<H)7]V
E[ECL<XUW,XU4GW8I(8PLQRM[c?TZeYfbB4W>fA94WbB<L[GVLdeY(^4I865U[\>
Uc3T;Jd_GLL#:aSM;GbZ62+7fG_K3B>=@\T[5bHZ;46-OaHQEc6fe5\?:HL+<ded
7AAf^F7LL99NJ<Dg5c8WII\-:J6JVY</KeXF2MEQa7dC05Ac.WCU7Y_OPDX.0CH[
^2O-[5ZdK1MPEY3<ANUVb_:N?@+98[?@GX1YSaF&RK8d@>b>E&gC8_:76O\1.8CB
Z1H#&O89a8cUFeNE<>GVOY[)#@1,/3>;J>KF8@_WCDWW]2XIAV#TYR@Q:Z?/(7\2
;KO2K5J>.AgD\HB2OIb(YX?P7e#V:HZ._AbHA.L]Qe[#G6EB)KBPRGdO)J)c09MV
?2&Wf-,5ggTZB,g;;c,S6KILP-bc:Z]aTS4eE-(_Ab:NCHUC]5C_IEHg>L3WP04d
^/T>9MX=0e[)O45c.d1RB4R>+PQP;>@V;=.^Z;GeMe=AT9@XAgd99g[EcPGEGNXV
5=&O.T0bW1D\4N5Bc5dC<+&(X0]\OMD2;P0[dRR;8ANXATc4\K&&cC=\SOGMFAQ[
??bQ_gF(MWUZg^ZERZcaP(E9d=e9N_(M@KX_ZQCf\,^BR4g@EUMb]\)5EcBW/R\5
/\N:M^eV/.>+I<<UA:bV^Y(RG,VPV+L(0#JBc;6C&abD51RV_=cG/9c#5a<)KA@5
3-?eMcP?S=Q_TELGVOGf^Z[03E#11FZQYQR]NG^WE=aA[O#)7.PBc-;5Zc#ATF)<
NQCdJ5C1JVKQIH^a_M)PY5TFM)QA:d3<4_GVa]GYY+Ib?JTdg#A86/R=E-N&ZB=e
F(B>S/(5=YPY>;0Z(Q:H67&b&<LEPVPI><[4/U99\9ffQAX9Fb4FU)^4+688B#dT
^Fc;E7gEQfCF.K0S+VZ8(R-E(dK#,/JR,4FRd32F#/b8&f<N)VaL&acNKEOK#;Ag
bMDPN+?fgV=A7SPU6KfdRf2^4R\8>B4fSdfg)a.3M]XG72XBd#ZD7++D+KJ.,aLS
,\MJQ>+EUcV=]@&VB/AIC>/3#_[<+DT348X\H.1MK:dXg/N)[7Cedc2a+>:Gc].U
HTT#9USf^Of9ANM1b@^L::Y:_L,NKbWQ+0EB6fL\]aKZ@A7KLZ?UIP:;E58PQW8O
a.8FTT^ZDJ^21BgCJR;WY@0dIf^T=)7U;0f^TR=TEW,ge#P?MY_Y9)KKFMAdMBXB
GLV?a,&\+D9(_+N>E^c/N&]-b(dY[a,+^[Eb[e0>[B?G_a[f2a)O<\ADe)Wd)fb3
C\;OYd9+deAX4E?\&?\]>;?7@@\2b#,5C\]F=b>SJ10PC#FZY2A>U))?==)4:cWD
b_T<((KWH9KU]-S0._HVY#:MI542I=[Y^-fL_6(]EM1.#R\RG>Dbb#I-a_+(9:?f
&faRP6XI=SQ[OB+ff?H+F7(^;J&-/7_:8<8F]DJLa&:IXH6L;+8b_GQ1Dd3a;@WS
T3eW]a>(Ce<4Ucc2Y;&A-:\QP-@\C=,&@@XRLS>3K>gJb=K,1W@dG[6\F9fI-FfZ
04c(0OA6#:2<5P1)?7FU,.ZKL&(PE]:-[bV+3E3UX2=bSX2]YfOH3f)=O&4S.:)U
O>,(@>>31LN-R(#3;4ETTF2P>VQY)BcC1M)aVFGLLXS@SXH&T]b1E>MYN6-M]&B.
+67&<P7dU<];Z6-a0#2Tec8,E14U_)YaA-U80CBA]6^g6@6LF4#P2)XX.Q;(a3\3
eI#,\IF&YF6:TMJDJROZ.a1e4TZYR9\8DRF]E;Z1XdVfWRQ6&fgSO4ag\7DI5+8D
X0VQIRHIQ>_9?XL2#LH.29+647Na3BR.,Z(A764\I;=U]5-5-AS.EQ<?Pd>cZPT<
g(LTVQIEF9<3b7-7bXY/(BL#OL=X&+P=:C4Z^)42EZC1Yaa1N>/8L[UTMSe)KZN&
\1[IJc,04>VcRAD>CX\GX->^F5MdGM(#8<M_3?-U(&U[a,c5Jg^E(@L?N&C9;Y;a
D-?O\d.80OIb8AFP22dI93E8\H46+E28+;7bMfPQZ^gUgS2f]H#L-EVG8X3I=I^3
));4>]H[0@AKV)&.Q&CME7<;6.NB[9IDJ0_g3MPDb6[P-#4BZ_CW;?[>fW7TdTNM
A_,Z0JO6fP1?2Kc8](Ke]Bg(.3RgRF\11)(XE&U]+]#ZW;dY=V#+M(b,IFB\c\[A
YDXR9TcY#,A;gF/d#OFY27gaK7-IcIGQG>f#SDNS=^@&+);CHQ@IAB?)XGD0IE<5
#8XLaISW4(LU0d(TV^R-.0d&[@]9g3ENcf_OTFLI2K@;CW=.R&@.?V_:@b@OZa[:
6SS9fNBIZ1f,7VI?ZL++4B;B/aYNCf-/F+A&E_5CVIKc/daD\CHL^MECI1BETE81
98?&T8=22aE^^a-Z<LTFbDY@?+6O?I[(,P4-<7OWT+9a,JY7GS<M9Ya(X&7DEg8#
6.\ea#JH)HCg[1I>]TXK=PC^Te_NL?LK<K:)F\Q<;b8C;37RX+&?gg]+/PbgPM0Z
E5g.)@5Y_&UZ]474d@UC9F1];@QVKYe1Y+f])gKNTfZ#0^HA/5IB=#C4;TM\R5A_
RXYQBJ--NML]W8A(B;E4R0_BU<>X5R15[bAb+Wa/e]Hb.W3:aG?W2\T1WcgIF).7
@F:UgX6Q.6R6cOWA/K?0aS.)RO/]VPKe;..P=ZJ(Q.77IccecLKXS\f=]2M#E=?P
c8cILY72f5-4SJPBe:AYL8N:_0H\N:c&LJ4JdCMbI(UC0+4.TSZSCd[.U2L((HY:
,9G_^E&b44AZKBZbEbLL[G=Q^()J;XQ2LZeW\[(;)cKPa41Y;3XGLB,Sf@FGQJ;G
(9+(Cde2/(-WfdF9aK<@I&T;1BP?HE\U@>-f](J^G4\)0M1HNT-b-?dda[[HfRQf
4]=L\]<M2,KcIUTSHbN3#f-/9.#>[J^&/67Q03Z&7e)Bd5J0Mb(/6TGO?=U;K^@^
>7J1M]IE)^H8dU?M>@/ZH<PLME>6[E9G8&.7Vfg/>0@K39KeZb:\L:XcT-^\c;E[
<Ie^40FYI2Vf;_[^+:+V=75gC([8aGHRAPIWB+<=A><7U-6RX35/P19a38[^CBe?
,eW0\EZ_XEX6fZ_W+^A,c@&7,bG,GOUbaV]+A^Y4Ig:;cYc,<F52>S]06JYL9QOU
,?cCf.I3GBSIe=0Zbe.DP,@K@[PAP2c#YM)Y5-4P+f4Y(.g=N6?G#JMHAAE6<U<X
&#AM>bZa-HUM-=-HY&.<_CBJ[S1Sc/)7\f4E,P[dBM6TDcgcf1>?@T5Bg+BP8OZ5
0Xfb)MfER8:1VQ&E#IN\=((U8UbdE]f)8GG?@J(_/L2EeKZP9^#FB-PHAJa4KU@S
MX<(Tg9e^LUD3E/dES[O9];a-4-NcJ,[QKP129g,4P9DR69,FA-YF-RA/ZK)Y\=O
QZC1&L:EJd/DN.+-c0<W;,0SV_=4ULP/Y.XI>SC::;\3RQK62/]9eEf#.4Dc5M\E
UQX#40Q;:LRI8NV?<@bWO)PF&)a-YYa[c:-3AJ;F?].d-,YRPd&37bG2I:E[V80&
SNWE.AD&Y@c?,Ie-,Hd6+V_P4&.d)H21bJEI.,\OAa\L0f<OS3>]2.GB?,FKAUNZ
gDASMP>(H<TWQ5JA3@[\2\B.7QB3Tf7I5+O74><S?5f6=]aeNF.AU;TYIMC&XQ\S
Z,3&7Cfa3/@+:Y=)ZSUS?[6H71R=-V)93HfcOLD1I<MJ@23DJ6bbg0d.2_>V3gMF
RH9DR9Zf,WRELbVF__C265AfJ368df:CRZ3=R[YXf1&(LeWY23D-MGEKe-)5[^^,
N)TF-THcU=T.B;I8bUe#_<0G>fO#T::9^g?,I&#(#0DP=G_W[BDg_Wf^eBB[H@>I
gTVMc]<0)RM2X1/BR/RQ>C1fg5F0ENM1_g<+S&D05MLW.-9)e;++dJZc5C(C.S=+
NQ)d(N7b0NDW]:EfQ2aCPe2<6EOR-Z-<JbY+QNQ[V/><W<Ke8,GOT9JYQQ&+10M6
/a(OJ/K1a6U1UYL3Q)@F[MOOUCUVbX[2E9Q?R6A_YG-IfSF:,H6.OOPM3=GBA#V@
[)+Bf<dbHPBR\Sc,OM)(\T/L.CcfY6:CNH?+e?LWbEUU_M.]P)JW)H(ad8)YCC(^
PRVD;5_/97fd>&S6>Ng+=CJE_T:T5Td7L4c-_K4TB+>NQU^fc^,Z-OX@Ja1Tea^c
5N+;841BI7T(XC:]&+#:f9^3PF<IW(GI^BOA+]DAB^&R=7/>94WC2E@SE=S&553D
A-,N[;,cg__@+LV:,2SECFCT8Q7baa_F?0g<\4Z,U--;Y1]e)EZWV:H,UX?9+a-Z
#VH?.J<+U7+?TaR4G[/)e+O6S_96YK@AN>?,YN?TPWdQI1ef;NFLG#ZHRQ(@N65T
fUdWNDU]@K+;OLRIJe7a#^05c\?7=2;BKbN/F/fO,>PJQ-EQNfebQZ,@^f.NgD>1
GGCKG=6X2gS7\21:@46CXKf9FBJI..U3/We#+Lee[^PT+H(I=PNfU4<BdcKbORK/
,LgR#a(E/2&>5YcKaH,4<<4-U>cO9gK956?J16@TVPER678V+(&^J?N&WM/fUFe4
>R#M9.FY2f5eDCVZ:,9/3_671,_b-4c^1RZ-b(.2L@XTaVUb9\:0\/YI3U04QZ10
@S&bI:AR@L/.-=PI/>]NYE2>OA1M-c+D6?-&\RQdRAU?#Y(#AgV]M^dRW@_)1eJ@
=]PcQ-PC67[B&:IFJ#V46MF7#\B#bXJXPg)[LY;gW,>[-K7NgJ_0T+Bd4\dMSaK1
O88C&E6F^U(,@T&I;eVdDe2H(J/g=03g,KB?.dLeQ-R)K)V&@DRNfZYUfZ\)3V7-
+._;A+(aN/b4WaEB>Q5f[WD45fXIFXFNc)3b4\#^7Ke3J&d#FKe@==b&6:2Y1:Z)
RBfM;_8KOONW=V1_.eWJeS,LB@465X;ZY:;-GMFE7\O+]d>SJ6UIR3,fP5>S(NER
(#14gB^5_LfG(8ZPbV,MTeU3+CA.JXgL(7@T]-A/Q4@\Y=#,:5KN@=cV?LL3e#KX
=a4XR)]51@DU0R9=AIZD=AQ<\2VL?ER^UJeb9VO5;BODgOFXF9#:2I:U9XO_@d38
/>+7G;CR/3d&:,D8Q89+#-C,7/\JO\PM@D[IETUf=Y8+-Q^=dL?4.;aC8#)bIBVf
IYM+JXBU(VeDH4YSIJXH&\6:_TH(9G9T&>[?572@aGf3;Q>4Y^<&3,#b6&^,EG+)
^Ob@O7?c4gV5V9bFe8>>ZSc5Q5HI<.H.2,&)>KFJRZ<f\8QT=;QB:WUN4ZM,M_XA
&ZBIaQ?SQ([a2NDH&XI>MZ1=Pb8aI+4@V5#P(>DR:11YH?cTV_YcV<6e>EEWY1[1
6X8<eGB7]D)3PN_MPJ;/T&?VgU?F<(e8:38^M#N-P-IE)]3=g?2M4X&L_]Q,2d</
R4?M.[L>O?DS^HZM8LU4O\LD+Qa4R+7OD#^MTXI::&f^OZGC7@#P:b4?&DJ>0N>C
[MIJ1X9#feFPO5U&#CTa=#?I5XIQ>#6NL8-AZ@CXU]^KJ2QTRId>f,BY0]\cbE#&
+&e^#7;S&DGSC#0C8XLU.]:MC46:EZYWVGe9YU[#Kge<dcgFG]V=&gd07=_T\Q\\
&6B+CcSfTc=^F9N<6X;5S,;U;ND4Bg,(R:#^3U_YUV\W]KY/aKVBcUV=O6+]W2S)
dfQ+L^XB6&4I+R1=Dd8gD8d?F@RFV68^g2(.-6ZZG_]P1E&OK=\X=6?La05Og\Bd
)/==cC>6O89&VBZYF,XYPWZ8^b>Eg#3+R734^a1Y>G=8?>E0M\-XLe\DdFg^_#CL
(YNMDU/0PV8U1_?\]2,AJ7-B3Ka.TH5+]J/U0K@A-6<M5)FCAZXeLGe-ZLeV7_VX
Y75-G[ODQKOU4]a/RLU\B7&UJQLMS-_PDF::L_^SN9[PTa14]Ug9Q\7cBP]>PgU>
83V]6IJ+DY>+J?GdGS:>I^2c#ET&5M2LL,LJ5>:AJ<=g\=F.W0CTKOQ;LRZJ1T&V
3+P>,]5Pe1AV^F^R7<d1+DT1)e3/8aCU=<.I0Kb][FcYL?94>^RJLe1d^^U;=Z3V
:&X#YB?P0#^#(NHINe,0\Hf1D8V/SOB)2@;2)XNOO/A&0:,PL+PRDVTXH>++fBZb
dXc7/\L+9R+U4_]JK7C??f:_SA)IJVe>@G9LV:K0]/>/>+B<R6AAR0\(#,WFDR=5
LEII.YYTc#IUSJ2=EH,&f,Ga[a7T3>28MWdb^>FO0dH[ZF&P/8]Z:5Qf-=[=F0e,
<c^Z5PNP?2XF86+/RV-&MF9+;?fJ<F[C.FD/+/-F.\_V]-,A@V)D]^1+A8.?_)G-
7Q:1?33HP<]ZP3DWg0^]/2Qf&UHP8Hf?d9&CY&I15)MS=X+&cg]\cbGdN2,RH(d:
VR1HFgfFcRU;A<HA7D@3e8#\/a4fXAOZ8c_--^6D80Hf-;77WJUS&T<:DXL1AG?+
-Xc9Vb;I2A-)abU_Ob&94ZO2]1Y7YZ3,<bCdb_\,1g^P:eU[<?W]A:A0ONE?,CdL
YX[Bd#NPd4-a]#(Cgc006&DOU4YPe<<RPLeTGDNNBfPfVKdGN/_a_0XY)TR;b#13
.L=1@ZH:C/,\AcBX(C5?Ned]T36Ng381^1c+[S;Q<<:dFPfUM,Me]TSbe=Ud/=R?
;4>05EF5(.DFNJGF;)4g>bS<129N)KPc4XL,GUU(E3<\,R=g]6Z02K35S37fX/?4
N#Y1]-2d]e4\cV:1L@>.8^99W1[ORUg^ZA47f9U0GIMf^V3g(+<Z\D,@(9&6#e5.
]..I#SZd6DNT4?+A4)RI]7JBVZ)1<LccJ_]>gYJV7&HM@>@Z>\@G;M6&)da)SXfU
(GDcc]>R[4CFR&OIO?8HELeP^9:I=UXSC_c\b=Z+KX90^TE<U[P3_R,gVVA4>(+8
e[FaJM011R>O+]E;d6HSZXWSP63#bSE#+4,Z)7DA73^gL6dE#)>]0-]8&[:dA>RM
GV,,B>_T]=9QAU,HUSK_J^2FI,e/L2Wf,QdS2_cV:eWSf1&8eFMC@cb&]W)W/_f/
I=V);I3Pe/dD1_,,BES]f24RDS38FcK=_7:\IO?[[E9FId^DIaUB5e\2&39?SLe)
DU)9:gD(YZY,I(/D]MTDS=KS?XL_ROWNHRWHJ@^;&d<E);:;D4:0.e<7e,;Xf?=U
WMI@)L?24_VYQM@O<:L9:<7Q@D#49OQ7.P>=Y6fNMCJF@KfdSW]#0Ab]0/QJdV1V
JZ=2@B^7@IL5F&7NU=@YF0.9gBC16@a#DX4?2/7E6\9&FcLF:((@HcQdffM]F+,M
:[P9B_e+)TI;(Z)c8AQc4:(0Y6+N2#;gA:T6-+3f@Y9RMVNg-\bFCD-IX.G)07U,
T>EOC[I7\N?&R-L+-5890K8Sb.-0c2cKQEEG_d\P-?O]?=PV6+0dGX.e<XCB?BO@
)T?O(OKaL1A<:45CN)#XV2)2O[ZRW>H-0_LQ9)0aC-LZLcb/_Ed712MJ)&1P4F1=
?PF5QJ]-^7AGBR_7.7Y^NeX5#;KZ[]<7Oca49A4<c?E?=XUEHG.SW@+UXO5<SS&+
&66E6Yf#6M9d)g91[IaO#[@61.geARV1]S0-Z>ec:f2LWN+,2RZVV3P#GG3feUEc
]UIT0M3+b,?L_K;Y)5+5LOGLU\@8MQC>)4]b#90-N?;@eI/M76UV-)<Y/W3bB5ZA
]MM<8)bF9D_FbZS+T_g0c_L_TY]/4<5M>=cSYO<GA]6d:+>H(4DV++cL/_?0af4+
PbYY1W^WSFZZKCb.dYZ:E<#0_09?I>;<,=L=E[<(^31#E;aeTI3d<W]M#6aF83UX
GWf5_AP3SK,LY)>PY.1LG1cYKATGG4bXMYIB8WO=^VWab1c1(g:3,d(2]aZH/TB7
LV^;&g1Jf&MY?>2V&#ODB^Of3CR2YHC>QMZFPXJ8,^P)Xb7(^#WKK4b<BM>=(;58
8(8L69PA@,g?EJC7YTeZX42E6RVCME_Ec1cVKEMCabMdW<60J1Oe?<\QBae)/.O0
4E\X1K-Q<([M-[&=Hg7&IRHVVZ+;HBPU5##,C1_2^\>=]<)NYWLOT+g088=F=cS]
/)HHb7\A;(AAMSc8V4U1<W<;T?-JWHN+XNX;NBJd;]JeW6/GPF\DDMC7T2:]ZMWH
1?Q&5.-&K[#L)F8+dS7EP#1^C@>).Ba<B+:(D;X9]+,JeCJa_\Q62L?S3BI3HPgJ
H)>:7]\.Cg-7cd)+G[c<Kg^6Z\8VR;2[aRDNKT2=2\CMHWMEaA]:_[F-9RSeM&+N
LUQ:#YSSV>23NL&-2F)LX9OE2XKVXEG-@Id/Z.T]A9Xd&7/D2J;DH_,8.^aM<ad_
a/PP@+=INX+#7=E2I/SVea6ESF,1&#<VD?=9Z?6.R),?>)5I6f63F^FdWAXJ.+5e
0D@([LU6G>OFP:1&C?I/g[F.1C=#;;4LFe0OK-ZcOL91K_KZ7RN+KBR=gU:JUQ36
S=af-cW87cbG1/9X0Jg>IbM4?IR3<VZb(d<f[Z1[DT@Q[MdF8PQ?.C5:DUE5#Y3:
\OGE9.^g6RV98g&?1(f_QbI&e:^6(9T]FF6XEQ:]\5IX&\0d6;7EbIKF;?8-E+>]
7eXDFZAHCN6S+9Z0N^9R_ZYK=X0&2])]f4<(MDC07=GN(]=9K]=UT.G:.4Y,[GD;
)346D8#MLOJFZR^OcUcHZ2(U,52,M_#^E5/G:3(dDJ?<LEGIV/3dNZd-.ZdB^0&@
O(N1C1g_8]f[HAg00Zg91>^]P_VNHRH^&.eW>L\J7QI&?L(AfNU5.O[5PgTQOU+X
8/KJP\FOZ^+]e7F5R/QZdTGc#EDFT6S2:B+ITAc<AZ0E+L5(@BaI9CLXf\JC=GcZ
@dC.ggVg:NCc:a.<CGfc.Hc,\2HFKN,XV9;c]5aECW&3fWa+=S04]b.I^CCF7658
=D(N-HL1XK/UPc_QM<(a1]P/bfUX&eS&6S[OT4AX^AL8+6]9bP.=WL79XD=^afZB
DMb4IUDSUABbX0<<&_\)4QcbI&c+1^A?#4?1>AO6g[OZ-/Hf0e99eJc,]_V&LUT@
>He8\)=K:&#aL/8e@>=@4V(e>WS6F\U@G@@\9)]8c00#WJL@L2_DgRTBMe7^g-,X
058Q3[S+W:__+2F?XN4KJ(acNZdJ^O220CQ@VH4^=0T>^,e^R]P[7e0##@NS]HK>
.K+&99OEW,b,1BU[DN2QNJIEBBcc6CSZETSXS5#[DRf\Rf8LSREd[D=?70(R&UIO
\Kb#\5,gdB6)B7G[[T9cY;cDdT(:?A51cRA3?a)bUTKBb9/DJHa\<WM6BYOW:B>2
28>:DQ+W=Ka^f?61HUW@/(8WTB2]\e0</<AU9bb;0M^YU.RZ8=TTMM5-TP?&9/5C
1K=S>ba@8C,;)R2M<4#dRH1[dZ<=LD<,]B83+Y\#;M;I\HY(e?KZ25#Ad8e&\45-
MA1Q,^eJH]4)BcW4TFR?T#-5S&KE.)@BeU#@XDJQR_F+<_K@Dg2@>.D(.1IBWD@L
=U_+E1B5Z&AY>f9PHT@)T<cRFg7b1NX3)c-#4^/+N1^>;768<]USAWX&IFTNO+#E
#PJd^-c4eXZ8C+7Q:eE:>R]Q;c2A)#7]ed/gF4D[.2b(CTR<LZW[We?P8+O]=&Q5
5b>EPA--ZgK;8e0O>H9BKDDe,Q8bPTS5PJEVgRE&>7O[G])1:Z[.7D(9<FFRM?S(
Kb(?O0;1^6G[7Ib?AV0-/fPH&\93S@H3:4Lb&AI?P2X7X7DJCCI>9&bMb./bC7T3
OH_;607X+BYEFNYIJ6OM&RaE7\ZST(R]d/8(eJ+,TQU[\+bC=2>:TGP05/^>F+Hc
ceW^/5I6;LC_R)cS9bODJP&WA;R-1\V^5>-UC3GZ?/<@GbLQL+Gc]c/0#3LM.KTE
?Ke:QgSI_DL?)ea4-bB,68b398@U).)865gY2C#6@.Z/LV=/8)HV<XT?B;-?5DJ&
W;ZdBZE?@>K0\09e:Q[^4PZO4[V9U)0(@^L-UP7A@?cfbIVU5ERE;>WZ4.P>[))-
8degeNGB/K\Kf,G:>C=8.&c\<[^aK.<DK^N2_cL3;7>K.DZ.4@1Z;/_BB<3.ABMf
P3[RF@V::)T^Ace3D[A4H9I_0Y/S/9:ZXP8CQ:M>8.X]()W0T[E-][>Q-]IM8=18
H6=d).V(1IW+NQGKJ?CM63aJcEWPC)2AJ5])7S;SPgP#W;+0TQ^EX:G;=I+.YSGB
5#4?R\dSX?gaJGXL4)C;I3Q5J(XN_;bJ)(a5RU7D6.BH+XKF,^K;=La8f=aVZ,T[
<RDb[f)]fS1X646QWaH:1a#]2;;.cYUCZ19(O9Ra,UHaKAf5@QfT61C]J8W_,@2W
AS-a76S,f<5X27/\FY,EE?PG/-Ma:KXd98P7gY?P[e&;CZUSM<2+_?T62#Y=]Dea
X?[YAdH2Ce6#5FK@YTa;N43E)2BAaVSN[KcI[<G<BaS+3CSYaL&#&9F(E:OV>O&T
HJ=IX+bGWU3?SR&1OQ8f()\.f54c>)X4NC<ZV(g^34b<OS@e7HRV^e9&NPDNcId7
?H(?&I3A-NUWLbca]3.-UAd.U]B1>Ida+2,<QV.]C&A@R,a9EKN89g1E09K-8)Mg
&e)(SP;8eQd,I<e9GE8<Wdc[,M?0_>R.-DH_]H5gBW,@PNb-b+@+)R\S4d,[<>W>
N+]Yg=,BcQ>[2Z_[#B0:\a7U7TP7Yf,,e:4@63F_c9>Z2#Ub82?-f4DT=^Hc(ZPW
P(g^J0I?bWMT7&[RZG6WgE+</8VILbM7H0DCWS6)&BUeJR.0,7_TY0(<=\/;@&T]
e\OBL\TT^DGe7/H)G8KE^RE::K?RI<Fc,M&MVOY8XI[cc<P#_\>W?6ZEScgU_3Z)
NOaP7<GeQPg?EdKQTCG5[gZPg+)Q>=(M[7KKcc?,9+XHPI_X@WI[b?b/914Q_EG#
/=98IX19>AKeM/dcBU]=TCVHa&AL/)]_@S42NDE+]C:X&W2ENC;bfg#ZO_DgLaSJ
-2JP&JY=J)ME26+:4&6MXOJ#,-HEH(_0+3EIH09?PRTEA[J<b4Z\L,ANT.SRER6:
D<1GeggfU3@KT_TdM#MK/^NDD_+_EgT0GO@5V@GV;/bX&K8#)LL6&J39fTEcTa0\
UM,]Tc+7cZ9VV,I^(;@HL0Rb3eQ,Q1C.=EHCD+/BSQC04;V-AE&)bKG:=d6H9)ca
,.3N;R8Gc;,,7IU/UQM?WSEY70#(Ta5Y>bD@f?M@IUNG+W/I=>/aFSQ-9[.A8+;A
7+/,ME8bWINL84Ad_#9/O]b&6<^;C,Y/IW1O9Vf0.Ub?1NFfH-IO:FZXGE-2O&JP
>TN76SOM;EH<RE2d4RD]NGU3(J<ecf:5Rb882+7#SfL&b4=>Y]EC)ROF+#^S_N=X
85)CIMZ#N0-SEIR_;/+^(^D8/^)Jd;I@3BRc1A/X48@a<T&5F2Q\BXD1N3CB^UI:
YWS-B_ZO2KM0WSfKUY:<LHgC,2C1D/5,(:#[fc8[H]F4bT>?<68?I?b?_X2BT]R_
dbBQ=X-S<S)KJOK+KDD3[]1f\I+?d:__K(R^:X3DQHSD,W?->5=_(64Y./b+eNeK
]Bf4#F,+^T48NW01c1\cVHW-[ba9RY0ef)]UCD-BIXH9?ES6.]61Q[4gM]VD(](=
bX77fV>W<H84Z(?V,:P\^)Q[d3N5AK?C..OZ1NIN&]:3Q4]3&Rb[?Oc0WY#,GC/Y
3WHcf9\N>C)_U?ZC&CYD>D4<ZeG]f>2Y#gI2TCZ>D>SKb64WJfR\f5?g3J6f66;P
K^K,U71/QB_(bSLGAX=P9bK5W=B^LW4)/><4W86(EIS2\UFC.^3BSQNJ>G)CPOaS
R[7_IdgRV#PgNVG[=I?PD,B7689Re9+7RUW(]e0M#?>_E5gM)YB#/H0K1^L;#7H&
W)VP?CU;)[1d:B#^SF/.^V)/a)cHV>&M+COXJ,.<d_Zf#\2]4H3EP;7LMD8&JSX_
c(U9)OINE-E)]6@IZY^:14GKDf5/SY[[:VU@@C)MfOS@QSg;fUg]?N+Z@H=cWe13
Ud/EXWTR2C^ae\B@;(c&bT^/)\/ggW3#/R4b4d]LY:D@B=HUMHML[,QM9-^3]J(]
G58@f)#?E@\b?<PEA+1+G9&fac9+&GF0JVW()4U4C>6OP6YR2([[RaN29HPdB5M2
_D&23YgJb,9G4\c;gf0,@d+_,__WB:PU\K:I8cC9VE\\SQF/[NB(I-^aTQI@OH3b
ccLV3W-NZ0E62GNDYK=.a>,XY@TCETbRQ\8+Z-X4E6[ee/@(JPaZ65_K0N,C,K1R
)5=\7\\)D\)=B?,&.IKYT:^O<6S.<WMB=CdU?ZT#X:TT,(S\BDBW_d^8KY9W5>(B
UKQ.>U,J@LSH,KHIL9SKL:Yba.7<MA<N0>+Kb5J-L8]gK&aVTUH@6U2ZZeeg2/d.
W>B,N)<_7F9QG8H0GV/.:-P;1.]CYH/7QfA\aRW060[a>>CDc3Y/#B.M/ON0+QV<
Q;P4L-Y6#^844L)@_a.NTaMB?<#e;:2&^FUb+6Mea@,SadPS(;fdGV+;1D:?/K(E
OF=3aOB.Ne:<-b^\VfC+OC<0P(&fefLCH^?;?W1\1C0I+2I;6d+@-5H>(<c1QDd)
<?V<7SaVH=3Ud2IE0>NT>F6T#3YdB2PfX[^Ja3.)Z80<[cIC0aFM8B45ZbT?--9<
,=M\a45G6&Ie2c=(,#Tg#[[T4YU</g(-NWXUd&]MSJ//.??f3VgVI;A[E[]P0ac9
]OT]FJ/\&87U4^4^g;MC4+_O^.A9+/:b8NaWB0&6cNg?+>KPBA-3Q-[&F2J&+U;P
GZ49\5WA58Z-UUBK)IRTRB[56>T@K\1W?,F@7L2O;/-N(;X3C\5_S^g.CN4WM=^O
);8-+13PJ&0WN<5bXPa(G+68.H#?K-[O,J<DA2O^_HN,]/dSeHDPY([&/:U>EN=L
3#b:_A5E1^MHOW;EQQ0.QVKNWa5=@8/=4PL(Za^\9Y4-1QD4)K7JQV0O_1ZUF^K(
06dO+Y]5L5K<\_S/\<8^B,D8BG:eb\f&)9MQOQ;eHSN#0O5P@D,>MefYCb.GB3BA
;/&/<=N>0eA^;g(EH>[e5:V]FM)Wc<2RAJ>Z\5fGFb?JZ?4<TIUK<3AbI#(b@_-6
80D>B==K2b?LfV[(Z@-R<>f9<a(BUDd-19g<?)=@(B-g8@?;]&?KdMEdM#]X9]_O
&2:=UWa802OHcbHb\+3PKQ6L_S1M2gZRN5T8I=C3H3OQg=Z?WZ^:Eb39-^-b+#g\
^5UY.4-NJ.fX01I6TLe&SNa7HR:^#1ad1Hc+M&R.#]R<8bC=-RQ-/(ZODP/]_Y_3
GKe-D+fE4O>TS7Zc?@fJ:;,D#@]Z+OSA)IT1)SfNR9<9M/&8<g:P7f1dRT0+RJLL
B7_=5GPI+>fO5)M(<+ML8eCC#I2P\,,L)>RTZ.H6^XFCV+e2HYR?^PS:7_XgT[SL
6K]G\W4<g[47f^#-MEAN.KNMZ=geSbT4<)eSW/>a+.&WUT1NIe[d3>_?>gDBI3?e
(WFRKO.S#1H+4\VM@T#^OM()9?IR1dOH/GNACLA?\AI/[H^,-_IR1TZOO#4-5=0D
\N^f36YN&@N:E?2ad\MU?,=V(Ub7[M-Y4De)_R7GHfD/Wc,B,+P05JP)]^@K;H\E
+_#[,gCPcOZF8=X,KVE5FII?6MBSb_7R=aTH>L6?C3(&PY@V5/]E/#gSD.d+E,(f
1P9>XP5.+N.6]E+IOa)GS<I@4GI,PabObIZ]:&W1(EYDU;gH&8@SM1DMJ@625T\@
fSXH#7?,&+<,6O0S2RcNX4)0d(9Z<IYE@B26?2((/E]I6-2G+#+H9SML4>UeQ2Z-
N],F@\:AaN/8].<.Z,1\CJMdPHcVR392.:=?.E<YGFYdDN1Y5+T#R.#a#P?N@EO2
O30<XXC&Q-a9-Ya<CHL?gH[LD-f=S-&L397WYM8S5K];TGQM7_:YYH>c=Yd&;eV3
_H_31e6SB^_(4,?YB53KQGH)1b0@3g_^]144I6/39ZAT4-S3H<Pdg8\gU^JCRc80
SE^1)0DN7MDG\ABebBR9XZ.(+61f(&9H]c@U(MPJ61Q9AAg7^C191]4LID2\8EC@
[USd_[X;9^M.8>S6QaU0>]d,0OCMgEXQfCQMD:8H1TE;^0:SQ7M)0WXVZc7Y9;U[
D#3Z:?16B#;L9ZeHOFSAC_@[(c2J85-(>5Q=A,dU9,LVbK(dQBS-^Q,MbA2D6Q_-
aJZL@H.^:b]A_@._.?fd=Ne_HM+Pg4J0:<6Z+(R2C@UCU#3A4#5XK)d/GN[(B=7-
@&:[cWg8H7DDGb?8I>X+^11+/ZNJeedC^I9dH8GG0)KY7IQU<HN6>d8IcT5&N1V3
g[GTBcN^A4I,)8@a^-fHAXcRCe&K_LA)KUHS0F8V,J<=1QQ:86Q59_gF/7SgY2VF
(TA4,UEC:.X)D&7IfG3VD3HKfR78<>N6IMJW2@?X?VGQBR-4N9QFY\:OB/Ga0\Mg
]MY#[3C1RU@C3?^L/D179OC9MJ:+/K07ZKE)5G_PI;4U6M1:<bZY=5#PHVH2:cU1
E2_Q1AU[e8H.]f5J;GO72bDY-E82)L#0bd6eNTd#ST?;V0S0^K7C3O5,=1g8gF2W
@9;Je9f6faK)J-EdO1/cS4]=KWH/+@c&M^O#LOZ@-P7ETa35g1b^7X[+7LW/a&XH
0;aHKZ4E<P^3\EC_I3KV]c>8SR6B&?9DUb:#6AM)Z7__,N<\L&XMbcUZ;fYd^)S6
BMdIBWJ4\PI:]NG3>,9F.)>3B@2-]#XSC[\XNVY@U8^:WAfBee]dfb]7DI0[)?=Y
LAUEAXB=0cSZ4?<M),,_.8WUB1>LN)gASN7_O^-6AV<+6T&W:XgJPd#KV;7K_La@
E/Ye#fP)dMaHGIN_8X_=2OJ;IT6/cSYN/eI:6];&\K@U9RLCQYafVGC^O]LSCF(\
2@a90WSHg9b@V34FEUZ:(1BUQ1/6TJ8G;Xc3Mb_e4a-?gLZ/?fY-fLR0;(Zd+..@
(],RY#8eDA1NK1bN.-R34?,:FA.U)V]KJTX5Q>[E;GdQMP8afHb,5PO#MOgT[F;T
&X[(.K>H?QUaQ?6P?_QH35?&X](]d]]acZ,U0H2Fa@&\fUSZZNRZP>_ZaXUA_59:
Cd.U<#B]gGEGSbeO8ZB.N&gI3J4&RNc9-K_IfE##L@;bCFUGK<Wb/<7bL3[0@&gK
ReR)V39/<3<;cd(HT.1)W+=C?VZ#71YXUc(W+C;BZf2B;X-^\d<;>Zf#6Va\<:7a
2Fd-5BK^;4SMA+PAP[a0DT\<A[+7KO/EJf\2<^T3.?_P:G507.VCDOd_-Lg^/,0V
GPMd>+BOg,T^;?.M\KaS4/686_,@C,+e/Sa#/K>2(>]aIR1=VJ#>A7?0-JAK&M,L
1eHA6DN#?d;]/>#7(QNbV=bP[Y5JaK1&ZdgCF2K[6<V/#2[J&_@Q8eAO)0B(3_b>
?@?Q@-43CP4KMU&O4N^6)L51H:2E6>f^e.aJ93^\,U9I):g(2IKZLFW#P+;HYfH<
.Ae_5YSJZP,42?K]bY+V1J]d1@Teg?eXaaRMD=Wg-GA_WB.8B[D>87=X6?LBI;De
[e>1#M;Z>D;0EeeO7JJ31-].74_BW=4d33Ff94E-DEg1A/Y>g0&;cY38+)GXVe(<
1cLEDe#c+:WNUEMB2/cSa<F\VW=Q(HPAFAYNb_ac6Yb62&C3DI2B>ZGPB72FWU5@
g]E?^aGAFZDNF:]5Z1a,4I6:D09?#=GGcT\ZJ+8-G?+]8&G5^RV#@8MS^Mb.<<>R
MD]E(g1SZe[\]1FM#I0a(-0/D^=-egF,OT7dLI/MN-0c);@gc9WRM6:bO(RWW-N/
.Eaf+4B0916<I3VMY6TfPSV_\;1&#(?:3aND@BC,<A4eEB4[\Zcg(]RA6@KL_DF1
Q_MYR]dUTKI^;3@LR>B7)LR]Yc2[#cERSC\DL\Y1BcP89bX=F)_//E?[0G3,O:Y@
;PV-ZR\4]aLR\JU-BdN&3=;(KY=gAg(C<?N2LUAfUDNI-))Qg.+]:]#4Y_QS->G2
/)J>@#Y8U9M1^AWRePHCFGV)9(O]A/MQ73+AgG07]\L((CP@->e).cWV-;Bf,ET\
6N<6-/_()29/]^]OTP/RXb0/-0^T3Z8GA/DIY7,>-Zf,H6DCAL9bP7C#aYMR^?/A
TJ4.KY&<_.;#V@OVEY<W+6L,8=@2PUAE1J#6[13W:R\NI=0C]QKEWf1;C8G#?bJQ
\T[FKdB<A\EANJZ8<9M@WPY8c8H#7VT(GcF?,;LKeG7Rf#(K(VKGR()QTaJQUG=8
J\?KYI[U6gL3^D[DT@#8@;1[:J09d\LS<7B7=/CfZMBJT2\XeJN],@+3H@:2a,JP
;aI=IK,-b#JG:#>]J>T:)MW>N77^8Tc8NJ9dcfV=EGM;MddQ;=DOaWaNVYW\=f.N
]bLRcdD2]F._EPG.@bJF8G0?:T]X:KTJRNO#Gb1/W;dOe#M6C0JNBSU8__LW9=6b
]UZgA97AHHaHG,M>1&b4F^6#3U8>H)5<X@GRC1@SaaY,+ADd=:=Q25W6BF2?b9(B
Uc;F>>,+.--[1DAY]YaH]ZG[&e=,:5LY1ge,[REQ/>d.d9BY;4+V6Q)WRYMSF,IA
[VR)AN1@b;K,S,#>UA]d^U.GAE.7c11C[2,:G^UbPX0g1X+6<B_+X8F1CDSOI0(W
VD++18X3BUZ=0UYETK/e>J^fN-8AJQ2IIY>>Pg^KKJ-1/6<2+4GQ6g_PJ4BZJHf7
<Wg#Y19fAS-#5LL.GdNNN2U>.^<d+cFM-K/R&)S7>TIUR;Q0NNb.7QbEK,Y&edJO
<M0J(HfD+gHT_.ZB@=<L\XDeN,62W-SC/AOfW?A=gc=@:X;.gT.S83JbEJc5.]X_
8/)8QS1(1FN\LZRON5&+e>-Y9\S0JfURDaJ@-H&229ePSA@<Q[O\#4VY(fW4g>GX
a0-Fb-B7)FQV^/8JM..>?c47E/eTK;0XZ5gAN#C7WYNePU:_DNFW,VVd^+<1aJNY
<GF^(H[4[L3\70e]T,LEKcg+==R<e0C\&K]V4],A27._6#a9Y-,GOdQ?_S0OHQ>X
\1^PL]b;L?JI5)FTWgMUC5H1OdKTM+4b@?&GJcV^HR<cIG_:f.b-2Z)>1b/OOR@Q
YUbYZOH#WMN;+;NP0VIb)aJ9g?U(E=HH;F#gPObe3Z)XJQLTC4Z?O,SY#>+gbB&a
THT#KAM0XbT7+0dHIQ0a[/0N].8]M6+.EBfB)5&6M2C#,72A\;+B<[Tf\I2APOaK
U)Y+ABERcC^4XaV2Ee^2)U/U7CcWF_Ge0QFd:WI0C4C6:7L=(3Z>G@E,-XCFHAd8
:YAV:=N+H7eM(?2d,I#C=fbN^7M5U/ObJH^aD/OG&SSLLbBVJ6;gB:[,Te^d65P)
/AG_P_0G)C1@UU2?/Y5?]=K-H.J@@f2->WJCLd90SXX.\,0E,7@0.&U?+JOeJJG)
N/KZ9X8dd;18[<aOf8ND]5OJfZc(TB.c>Ta.A_^aJ1Qa5R157adQXPfJ</WX2HSe
)KFO8YJA@T3?MTS^/(?E,&:e(I<HI.QMO)5A5bZ_20KL6#N]>ND>#0aFGLc#:BE+
H_EEd)3)fd=ZYXdQ=N8+NE].gcF;+/:QH0<W#^X\IIEQ##Oc8ZfT8UafGY4NJ(+7
\8DSN9@RHYUL\5ZdL<:^Ga&-0[[MReFf,I+?OAD/LG4@P#+#ZZD#T8^\Xc\:_C&K
W60dbVAEM^1>\2P9XN8&5YfQ5>+9\_,.9P(LAMR/(b1XV,CTV5)b[IWEI^VDFdbf
&Gbg.X&9U]IYa?NIf2dQE(:=)aP@&/Ge:X)IO7^))a2c.CF7fN+^IRNZ&-\;S,/G
9=H+O-&/M;fOVEB4R?(?MT5N1(;/PPf^ZDIT4Qe<K]&=_1J&HQ=3c&U>c^VN2ZAI
J3=L)M.^^SUL6=)6];1^OF_9S-]46XF1#Z@P:XeW@Q+DSaHH:(GZ;1?ZG4TO.Leg
\1FO8[fa\/@gV(W;fLVcg?(17(4>U.eEe^;6TR5V86I/7JE/ec<IHU=,bfKQe2[Q
;KKg0.6WI9NE&VD>@cWNG1HLf>MeF+0Q=(5X93AC8?+ZKNBBLKQ=CN,\FbLXSSF#
cGb&cd[H46,95>0M.(+Pg<C[/W.^OB3NOEU0g9O=+8WN,&F#2gI&G(@)4.aI^F7-
O/3cIbGVV899aGS>Kf^b<)07TcgYHJFJ+R.gWM/FJg]09[c&>_KbbX:3J&;EV=?^
8=P.>.5(Z:e&M^\=-@K563@dM@&d4@\?5Q[A1?#CM<Z/aUP7^.JaecfM7..2TRPe
=66S(3dI/fLRT:+)[F&CcT2HWV&Q/K+)QLKM6)g&02W3(00^VVW\=/D?M3;W@&#E
Sd;0Z_DfX^-aQ1X59)F]@FPC8Q@@g;4&#L>O;NQd1SB&aGM8V2O8LbG&<g:V(LSI
A>EQ=fd)]WZd\MJ#+C)Z3(K2g2?;-W\<YTGM.c4I;bW9FcP1U5+U>0SYHHa5?S^(
)Rf,XfKHLQHH^^bHG&.9X\TE@]14^AWd4#FfE&X_HgYLSYTW\_1GR-MK0,[7M?LZ
RAL(5CE)^OQSGM)Q@0HcU&HRFFY04S3<OR0AWMa;bXY[N0e3;U(&T_M(?W^EI?cL
:f52d0A[AeQQ(<GZM#YT79+_&+1K^1fQSWGZ?-@RD/+6J1<g<G)YET_K5\+//EC7
]HKEHdVU<)-(a528TV6W&F@W3ND_)TBJa&Va1b7<L3HH;3a+#d7_g,@f07RcY+C#
UF)826.(fgb_#eb^?.:9P/e3NY(geK2V&.a7Z5K5EI=?506Ugg@SXeFcZKE._;W0
M.S.V-Y\@(^5R9cT0Of2#OTeSA?^@8)gVE[.Sb6\M8/,G?)WKU+b:FDTP^eWUPJ=
=\c1[:)a(9&H#YD<59=RITUK9;Q=a-VH+4X+g[TfQ\JP^b-&f#H=UIMNc<=C3/Z9
(8-H3?Xf&9C^._f]g9/3=/=LMI)<O1AHS6g>FAX8gJ0dSa5[76-4&ecSWGR#=K-4
3?_F>Le^A?:TRQ#73gfNXOQedB^0[aeQ.O([e3TJ#C#CR-3RXZE1W<VfYNM3[K9a
=P^GVB-Ng7XM^DgC@8RZE>T.W^ZcO6,,[&@+gU7-<N76VQ?,L94KUa6#cX9/.;AZ
@A//6,A[-9OaZ@J,P6YO>EJTBX[;LZC54?[dFKSPUQ>M?QH/aGf7;Z3WVN02DW.8
.O#2)JP7=0OP:XVDL<J3(+[S]f)ULY,Gc9\-28)31;\L[5ZRYd-Aa@]Xb2+HdBUe
Z2#W,19(]P=7AXg1+[;&E:Ug9F0RR#=:?J^Wb3C>.1LeTf74AAN(S+b[-M[W[c4B
T0VXIP[=3#cTCaVL.VXdcfJI3;#):R7d/>1#a8&DUGSLG@U3SF/=H84M4_b<3ROf
d[OGTS[4J/][2#dZP5(NZVNFJUIf_Q0KSKIR->XY5JdA@O4df1U)LPWBCAX0Rd5>
IB;5+#RW[\77BE5I#GH<O/A>3I4AI(Q:R92G6]d]_L:?B1dWY,.WR_)YOba\VPI3
a>JJYGeR<_5FS<<SeVVRE@5?A=0>NMG.T.DSJ+U?)_U,.95)g_05P#OaQgE3cF>S
aG2d<5c8Fc##;=7LI7<VIF4a?)3MZ;+LNHcDJ6@N;]&YW3/9]WD^VE/S^472MPcc
Y?S#G:_<Wc3F8TO\beIg1SfeL<NQ#F3X6L1WU+(;VO\A?->L9__((3@=LeIAD])X
d@4=5Udb6A13XQ2E8CF/;/RUbJc=Ve7d;g-;9F,;045HE-LBLY/?1Wf&G2D.D_1>
(Za@6?<@g.<gB(FgFa)_C((KOa&_Rd,N4Z=+Y9HUBP-C9D4I8=4ZI,T6C0g(f+[^
^<X@fTL-2L>7][DSI3Y?:/H;\bIR3THPM:VB3GLKT=&b4EW1;6G\;4e:)Ke5KVed
J&)@&O]0F;#26AB,a7(Y(HE6@UWec8L[76@&X(2ZeGKV+UNF]6-)e[.g2f5B/6J@
5[GgEc^OMO_/0[V/4c8U)/P3^c=;.]HL+4A=4d9@b]<N-EC=V?eS_F,g6F2a[3[]
5\TK]9:b3N[5d.K]V2\C-R1,25BU7C]#5/#BI_a&)#L?PCVb\QAEZ+6U0>>b^L0(
[g=:RN:B4=R(gQcWEK<H35fUR\VXC65J/<.f^G:]./MX,\BAeQSW=&8e>Wd^8EFM
CH5+Ve:9BReW&XF\C6SfP7&V[Y#fF8Yb><1ACA6:.Z4OBS+D/Z/:--F^(7/8<+@7
7)7eU^>[;FDED]1IfN+QNI//C\J53OPa8;5&02-5CMQ.UP?\_VN3\2fb8QET9IXB
2?A5OT5I7;dSW\bC0>;8:/84+If.SI+>^\M+52<=5f0U@,6G(]JS?CcPV1:C)B4I
=7^?d9^6^11;#7VU?1-836XQ0B^2U\EHR7C87-W-5:fXPaBM\#@eLZ=/\+\d4=&]
(5-dI)2GQYP#,ceI^Y1?Q[R(U0>4,S-PI#/1>UgQI_7S_EHbLX#8+MLG>^8N<?+#
H<@WXQZBWQ9eaT]NDH_IH,[a23AaE,5O))gKb#SSD;)fVSU[>AX5MY,LVQY[?X^6
Ve<gZNX(8M.50#/0OR+L1EgHcM?LA:>1ZV/2O]H:?ZbG4g+3O2/KU\bbT66_NL0>
M?_B@0V>@&9CEGQcO[P2GROGGgE,J8KE^>>DYF&ZVXZ3/a]V,52:-e^JMc?X:eb<
X,KE2;KFD9<GOD<JCGfIQM+#,EP@[EO5:E7\6R0C/9,<gBB^X7&T35H9TdMB_M/2
5?56F::dFDM1.BT<G5&A>P^&4X1][&@9&c[4J@UFD^9T1\U7YdN>_GP<F/#S]Y;@
[3@,QW][)O#.).[+f:6S5bd^QWO[RLZdT#B#K/ZdMdK^<CX?A<QOHd,CG:U?0\QB
?X7&ZWaG^8I>7-Q.\2J?O/dRQ.M(C:_^1I@1:\c\F4XS:E(@)d25.U?TJB]eY3OR
@-[I:_8Z?F?H:2]ZE9K0_.C\8.VNX>TA^U+08G9X^PAB@:BA.=ABSQE?f044-Q)4
1_,-9N3LU1?gI_N483F1OVWIB^WSf+REP5\=3JFe]##Q5YNLW.(GZ).g\_JL-(U7
:#=QT02Jc7/[+cTI038a:03.)>>9SgcB7@CI;/1/.V-F+V)&SPIFIa6Z<.>BLAN?
GJI8+UE8FVS#e(09.M6VQLd,#0QK=f9b)(<d9Y\ZM;b>1d22(P>--<:YO:7I58L6
XNG1T9OMOO:G09+T-,#8(1:5=<[A5cH)^G@[#<8);^N,N)6L9ZMROF]?\J]AOF]P
JeRY6eb3:6,61b>[/?4O]&E)Q5?=P@aS1HJH<_>]D:)):,4+:/2(gKG<YI30H\CQ
QSOHcS6(gFRUc1f;(=aE2#,[YeUEbCE(c]E1\cH(9<b)b#=)\XdUEM[&4D359<19
ON4[)-I7.&L<^-WG,Odb^fYK2V&^O]/HA<cQ<NCdWZDX&@8L&FPfW1=#]RHI0PAR
>D9FWfL,)_<Xe>)H-(B^OABLNC2A;<=PO2<3GQSDb;[U?YP=e3WD)Z6,1._Oe0.;
ALZ</]3TVP&PRZ^#(FPAIKf+L6F]GR\.\\MWL>Y#6I7W.]EMP(Ja3:LN,R<2f]Oc
/e?&QK&bc:Acg-aZRCCE]e_(:4g<eP@a@<VY1]YTP0YCI)J.JY_G4E&0JY\R1TP]
/ERd:LJIO4d2PYgaE&)_D@F&N=BPHBd5f.H6;/>&#VZHA5fXLc@QE/>6,V1BBg#B
aC.WA/W;&&1Z:S4^\&/9^YdPAfZT,:,UKJ(,\>E7FbLZQVUaaQb1O+VR9>NJ]LV,
29UdB,7Y2U&V?P9f[>dgHY75:Y)F_Ja7M5N^Va3H0UgfR\G7#2>;-cJ7I,RA<^PD
#.f/^;N26R-NYVeJ[QIA6T<WKOg8TJ:&T9CZX?>FTT)NO;H9I>#@QfN#J^][:..&
HP8dFe&2V)[U>WL24<.S^>CV&M[5U2f1&B:9Q4>A^WN[U.#=]4V3EFBa4@6U]N/9
905NHN@])I.O(NA/4a]@9YWXbReYYP_/NZ(8).2FeE2_?c,Sb-R.-5BEC,3G.V<-
f>1FX?;4IC=R.-3^SA3B8b^K+W-?N.I_9XO&Kb^bg;=6PgMBd2bbP?45DA8d/dc,
D+:af7I8YY(LXY5W.)9a8-e.G)=MOOI_B7Pf>9\C<;V?GA.?;KBGMc,CR^7RMf&-
)W;I@22WVXM5H<T#=;<4+OTOeP#=Y[W8(\R/.f5Zba\&FZI.gYFS98CF30#]VF(5
Qd]W_#@dT.-,J+J#W>E#_KA@/KNI?GF,WJL]PFGeFK)E.a15.K\J6;G@,>?>H>+0
W?S&GXb:;CL0&DUb+b3_&3a^U3^DQW@SaO[I.W&[1F2U(>W^8)U(Uec0>S?63WH.
7C#GT8779W[7RP]HH0FBVgQOIBZ;>+L9N3)L)ab,Z&;4QUMb6<^b0F-1TQ95dFJ<
e])W;SbJX#Dc.b\.?FJ+U>W&7QAE<&@/4>@8gED9-WBG/3,gR;AbY\Z\@F5.e+>@
(O:;6ANJ^KU<ARcea2Xa#]B4&^^CB=@@0I9HNGON9HC>KHg=\5>(\(gC:9RJX1He
+D6]2ZeeW1,K7fN]7YNTDc-TFB-0=b&YX7+#^B&>Oe/=Y#\;0@Dg,7-H)RfFBO+C
K[IH86AL<OBD46K&8XQHd2V.X123PBB&59_5ff9-b^T@VJLZ.adC]&7-d8:e2+IK
09RRE2ETV&AG\EL<,WV\_3G^L-XggRJAe3aOVd#9b1K4_SAGP,]1f&bXgC/g]#I=
:C#A?0=AS#RUA4d[7C)bbg7]cB&BF\d/]FJZPZ,,9WNC6&T?dALN+W#/5W_Y7@S8
Y/gBEAG8\Q=?Ld#WF=+_6(9AUQ(gH:R=WIOb?S;11FO,C\MS+&[>;2_9H]\V&K?E
W0-VT0I(/B@29.:gB6_4afS=&Z+/gUM81?MX43YN<+MC98G98Fg9+T48_+cfLJeZ
KXF2d&Z_d2<H2Zc\/WKPMd#B.)ab6=>-1HYLVO.+\?_fB7+#++]M+270bO6^=06#
-ZD@EZE1.78Y=_+fb;.aUFAJFWY+V<(.C)RKVX]:SgUd=P\9HOGe=1LJeT?)F:@Q
#N=]>M9IYN4F=.5&K0C&3^POQDC0&H&Pd)6[INYWD594,da;[ZBJ\,QL/)U\;[T/
1EZ7dSK<R]</V<1XV)=)NC3Gf+O/1[X>=CZ).e\HI2b(;0gDM518/JDaF=+3[H3d
?[ST.1D896bd.c#5KZd-3[T.I&=J8.GG7M0Vgc\E10(+5Pg4-G]V)A4I@#;JH^[3
5cE(([YKEIB]2X0PQB^;)-ff-ZF7JACQ4_\<84AI3U?NZ,;caPT+We3+:E]d/7(J
XNg4NAA[)R;?Eb:?6(d](HKAJ]Z?Zg1L8TQ&GW6V-#)RJ#NbAX<WV1ZJ@KXc8?SD
fG]+FWY]gXCf0X2UPX_9=92\@+:.c_G&&UcNE2;]bQe_VB^IMNf&;8bXY@<ESE5=
+K<1\3G_U,Z1XQa)gLO<eQ4b,/1AX>3XG),?;],9AHK;dbCS56M(SIL2Sgg+X4BM
8-X7&MD/d-Mb3T0^dS9+35)BXZF?6G8;+K1We<W2HOTbJ;Kg>6BBdZ(Hb9[02e\3
Y:G@AK]C9<5E1RS/+H<4/a;^0+2-PeML6(ICc+NC+OT:6&G<8JLNge6O:;XYA<^a
G)BEe#YQH2\e.&&aU\)ES>O<M2\Sc8E_P=;A0:QSCLY.&90+,f1c1FW-^@0),JLQ
S7./0;Yb]@H(g>3)a#FMe0K]V,;M1G<3#4c.+-aSC_KN-eJ+M1c&Yg@<F(W=Y#>1
Z^78C5c8L<:FZQX6288b3=&a&S2:4g<TR+IPQSGC,;\.@3Me-2B_TD+0ZKH04B0f
W<42/JGa5VeA:U2LEVN+-KE)-e2UJ8d@U-WBI2HEWHCg#.\BeaRODOeE^(X:Y-5]
U7+&c=2@=QA;]G)D#.<&Y.@2.)J.7&Z/PXR<?^,TXaR>gC4cS>G&-FaEYDK;.,eW
)4Bfg=dOMTJSFMg;D[--OUBga^REY+&dC[D<=C0edd#QH\R.fdOT>JT2LB5dbJ6V
[a<R,@+[_?OaN2.[J[O/PI=WcMGE87-&+L49F9Ba;H<#]-cXNO@()E+M^:@HZ;a^
]]2bX]WUW<P28N.SQ\7+]#2RO^/M1NK/KJ3E@+_0P\3G+fFBJ^cB)-@U#bU.D3(+
6N#:=fXT?XdUK6+:0H5W>GS]T.b8a6^Xa--^F/0=/_B]I>VdK9<75;@[J8NC](TA
K.I.(,fbbI1ge0gDSZ9aG(,5,@L(96Db;4Mc=W]DP(VE[UD(0AWAHO;[,FX=@&DZ
b:>,1P8?<2I\Bg]+Ob?cBG]CURN^^^<SO8ZA@D2edTH5QR/289H:Q_gI._/+PPA>
VA3PeN+J?^Bd[Q/:_+E<,D>O,6U&:KL/+>]T5H4V/>>:2=_Cg:6BLQ\^T3/6LQ4M
?S@[c1CeM-O)JX<P:0&MHK+UG5Q>IX-WPH-L658J_fHR06cYg2[JDDY&XCf6D6]c
Ng]=QY(HY0?,8[&)#1Y:^F[W2Fe;>Z+GW;(\LQJ3(PG^F6HPAU^#]:F0AFHUWUE+
(TQ]U/=Ie-fOF2R(1E5/D;c+^T,OB).<<G/(3-9HEdG-(^_&d@gA#AEXGf[Q^dJ2
d_AG\:6FHCdba#3V9d[[CHST7:SK\W_,_3c>EgDe[NMZ_[_&?)=&#\8>Z#6F]<)R
:<DIg-Z?^KRLd_^/\R-JV;F0gG2Z(&Z?9G-0OE+a026G:8.#+g@SaAHUb13g^Pd,
6f@3R(bHPBP6KPZNEcRGYAcH6A4e#(YX:J0.8_VA?&bb2de=-,V/4Tg70L6O(&A<
M@aD?dAD#JV;E#88R<92_YISL]-f-c^7G8GB)?,&Ie8ODa]TOPM=D?fO_Xg9gX97
7DQ.eZ[?U[dZ>YS&8;2-T@)5/HHRJDd(?6=Xa)b11RcP7VSKVP4;B.8_U6^Z)CW]
FE3D_C:GD&5@1OV1TB]X)\_(g,F<g]#-\Y_ZZ]e#G/8Ye_3a^6&-P^_fAIcZ@<(]
KCA/);e4,5aUW-3Qgg\)1cZ9MYY23<-8cF>IC-;=[FV5TRb2K(WD-af;8@A9&]H6
QC4X[<^1LQ1F@MPRB^_]>]RVHTaM#gV9@ECBF:6B5dPfc[/CbA66R_&T26--AdbO
=gS<:.V-7TE_<S[:]-Q;^A,FcTQ@Cc:B52_Mf75,<-#8;1g9;[3d?YX<JW;)U3].
/4R-2efFJ<O_:,J5I&+F^RA0LK[,:WLY(=X)QOMP.9RG\YUL:\R1IXfF=RT4?SK#
458_^Nb2R\/U8>V_]df8cYP.<O:.8_Kb934H2_I0\[:GQ6\@5MV^]b9:a;=9R4&Y
]ZeYX.=5:-agg>.30P-5>gb.-bEV>_0RH,7H@R,O6UfRdfe(4OM(K8RD2,,24;gA
B@g_CB:VQX\8g[afgA(0=3f7)gV?IL&e#(</YN_>[GYBXMcMJ@aa7>?\R\Pe1cGF
,]?U.V1(E?34W0KB:6BVM89P?&\[\,CNe(0I)B&\dGfBWJCQ/=;@dI/U3<7OTeUH
bKC^a:L^79-X?4,8=.LeMM[ZZ[Dc\_^+^R:X)\JTTV]>85dgQ-fMY]@/B:E5K<eV
?7Nc#\GW4CA01&VB>CWYYeNFH4g,6Z+7fC<7C@YZHPb0/;a(M3X:e7=0YLI7Uf;@
HJ2Eg1?,V[-?@CA>+fK5Vg4N1)cFEZNSdDODEe)F#39VV>NdMOdaTR0eZ74RO[86
SFIF_@+eS^O<BaXO3agT#@Z:=D-X?S#_O2I^G01T<2:(EF9.6+UKe1(:;S)NMW[J
f9BL#&&0-36C3CM07aV@+FFe[]J]TWB7]b-(QbYKTE_I1LHgAQ6I]+]0bU9/JK57
2EX.6JLIWbd=Z.4)g>>Q:105&N,+2)],-1b=;X=[e_X:9_ffTF0#5+dH_@E_]A>/
ULO?G:-&[)GSC=D,c-f,42dQV@fOc:U2D0eOL&XZ_<-RQ_G1:88=2(^]7+_)L_L.
M>b2CBJg:B[Y/7-4G1_WQ1\0H04c)\LGYW8^fNcT4G+]07\[UB_gPCf.<6;MR9_H
P)YcFPd4b67P=3MFMgZUggA0V0^8fTU;PP/-7]+Z]HQOX8GE,Z,9&/>\+7K+0+;[
G-:C/>1GOA##)1#YIW+F^:fX^fGYFW?#2dOHa8UTPK>Ng#b[+H8f80V#PR9&UO6@
V9d,@cK435@XU#K@H>^W7E0979CG(2I^;JAV-W.^Z.OJ]8:B9TH7<H=&6c8IC<DZ
57\QBaY8HLH+<JZ_BD)[0KA.)CD]1R;5Ng0]O<[\FWBY/QXW9fW1>PJ+>^OP>R)G
gS]9<4LaX0+4&fZa<8Kb7EK.(]_8PO_SFNg#gR1f4MB_e&TA7#&6?b)\eD?EPQ3W
<,=J5a6I>OP6Y(=5f.]eIJ1:G,-YL_0eFg<.XfeK,5c\PRH>N2,?VYYUFZVRcP&P
T(<RfY.H4PeUP.T>VNfHMe;FVDJ-09BUPYbZ+T]&OAYP;cEIV[fYK@(J;,JL?b[-
?a&95=^1;bbc+6T<aO99MH6<.M<4dM&+#aa\YJe9&^?U0FHN+=A/SR5E1UJ#1=8A
U6WcAG2ZffCF,FP=C9THX@=Ke):C+8C1JK_.UN:5->E)NZNVNUVS9\QYFU=Ib,8M
ZCS@#JY:#Y)DbCMcATgY8902(VYgK/b-/9[e@1UHOTVfHfI(8D:a1R999+dYNY/(
62M0K(CDd9OLL1T^W<3:2GG#]fC9M\aVC.Z7AV[7Lb[ZR(f1FM,WK&_b_ZU4]+9O
[#321]#Ef5E>)-YX,84OE^H&B_Rg=_..gWAYd71=X6??LG^c,NfKR)Zgg06e5.1Y
P:]2LT(]eI;R4(4/c<P@#E4RU.Ub#)>Vc<[+UO9>b3Y@W.RMJR<;ORAb]?QYK@8V
eQF6eL.J@.e_Pc[JYK#TB@NVJ:Z;QNV>YWS2aFNDdM)/0Kf;=E/9:19D]fQR2=+7
aA[^/Z8dV0H57g\KI:FF8HZZ[@;\MF;A5PRc7b8P\@B^XRE_6).Jg3IG1G3\.bTd
?a\Bf_ARSR>1GUgfcQe#P^4WO4R74#g[+U;:CY,P?QVN_7dU/\[0X\VHA)fXRR-\
cTbd)_D4@;R8?a91_>Sf/Jgd6OR.e7G+KJ:TSZ?fLg+DU8CeV_>U>PC@&T2M1aEF
>.)d@FdDE+LBOeQX6#UTK5U-Y[,BRf[(b5N5BD;ZQ.(?U>Mb5VBGI])X8MRVAXJD
GHIO77-)(/^3A;B0L)>G1--Q,5P\K=\EO909NR8b>N>b\\T__f4FT8f5ES&&:LR_
6BKP-XWe^5Y/(;U=Z1bUY(Kab:/#c?9dOL.cQ:Ia,F4.-168]1OWDRGdV\75[H&G
9?_/WIHZ:PS6I+CE6Z::C]2d#0\1dJ=,(c7Z8e>?47V.K944^560L7O6X+fDeX&B
@W;UY8BK4CM][P.&L5c;[PTQ08JYa(1N4F[Zad\]7-KR?ZF;NC)/1OUB(KD=F<@\
<M-0LNUFSKUNV;>ObLg2W0^=MAC.[(Z[PeM6Dc5DT4\E5VAV[FE&>f]&L2-6>ec@
1XEg8FHe.&8KBe[H^YF8#_Qb+2BAE40(:1VF6;_g]bU>f6#R[EQ4(DD5,aeBO0,@
0a9?Z3&4ZR[(d8e?A#HXKIdZB\cQE0fCLAdDKF(:8Z&G58Z-.+=W;0Z3eHA7JgA2
.A[eMK0M\@-<K:X:^V]OHK<-F9CQE=&WfS5O.(2@?SN7L6W6bdZ;YC.M-bYBI-ZV
R^]:dLC-2DC.(HWG=<eQ8Ag0^G=b7#PdS@GP+04H&U:AP-]_0LAc>G@gEI.5+aca
S[Y0RP\3)\S_X3-?IG&SZC>QLf;e>W,C^MDTF7)XNW]LNF(8[;_E83Vc0TURNT.P
9XAKG>JE4U5.4UNQA0Q+\)^[HEQbW+A[T;-J_Z?DMLZH[,;@FHCF)PV;Y3U-]He[
7MZZ9OQd?SS4eCBQXBO9g-\CXV32RV>MKK<[3^S?W@5:M]Uge)<N]X.Ef=FP#[e^
+VJ4^LG2;f]LdS7TbJV>\HP?_g77M\[Q@.RFHT+gP/QNT?=b<O(AJBZbK7IHZZNc
f+K#\5F1e8_KNF#?b]FEZ(<I((RbO7.cPKKXKF>7H5\J?d)aEW;342&V=\6.d(JK
aXc4/4g+d_(Z[BFD.Hegb:g;_&dWIUW0WEQ9\/?U<F4/YCID=^5UfJ?<RB6N\Zg6
[?:AXfJ<8YAOT2SI1NPQ.5IZ&>ca-M8<=?;Ag6.26>c#cMY@bDB_C0:eGUMB6(/]
PDZdNH:#D.2?S;=.@feKK&]Od\QW3AK;0/c@<9V36Z0a#f.f\VTOQ;&Q3?.QI6E:
^(^8H/747AT0AZE@.dObHU@PXIJ:=T]^:b&H:-a7QE,O__J#ZU?3M-ga4d>_HOM(
?YZ1Sf1W)W+?BCUBF=2,9g:10,3C+eV22LIbQHZ:ESF#J1cYIXWO,;KN7;AL=0-c
?#-?J(eD__4Y>g8TabNXO<E<9a_e.HZ2>c9Ya-b6PK.3.(>)4G9T_)550(.ec42F
O:7SR0c]Cg3BBb(.6+LM5UFU7,:-BWEeX>Fb^4?[a6)cJ[C)Ua5+FWeY_8-OW3?P
0S\CC:3)HQX>AK6>JVcELIDe/?PZcEFJ_>cZFV,4B+b&Tf4I25e^Q]L,>-6IG@;-
+[[>Qb8;Z?BK9(Lc83bBG\_.4E),@LOLP<H]7<bE1C\PD(_@6I=1B<&G-CV5_)LE
g:I62#0;YJQfbH2QTP3fGQUONDS2=;):fWQY\,#;e;d3)DA_Ag:FWMQ;T,7NcFGO
8=.MVfDR-0(G_7+(A8-V:+5[;W3MKFBd)a]#32gcLVVKI.K5##=A@XbX;NZDP[+2
(d+Af;OT\:Y9YO<,C_BB?/=_S4W],[E<:4Z>P2\QeAIKB<O_Q1<^KVQ^V)FQ6NH.
H1?,]dR@Bc8fV&cK/CLSC/#+]3V,_YTU.W+A#d@Q)VZdaQ?R+YHAJS+9Db\ZC-XE
CM1f@PK4[G>g?8df:ZI-:N2_B=ITg<]+3#IC/b_Z\Mc9Q:LJ#cW4Ka?.611U1<NG
L0gYFDDWAg<;Y9F-R^f^+&)J#)[T15W/AMfL=CZAT3#SHDM#(E?.E;4Q8J\U?f6;
HaGL:.)dM29=EaEH?XO036[C9J+8LV]X<&6N87-6Q3=gbaf/I[=Bf@eQE:WcH2^F
>+X_b5K@gOOO[bGT8,6+J]-Ya94Df(N./G4LDbb+bLOH]]:H(1MCONI7#YN7P/d=
g3BIYG_MR5YXIG]Za\9Z@]+6CAJb#?a&7:+B+.e2OJ0Q61O4[EV-@)IX&aWaCAS;
&JC^SMM>ZP1^6L_V<P2_3WYRXaSR>RWY:^0W2]Ue[V>^O>TG5Q)PDVG\EEg9&=H3
<)M.KS2-#5]D6d;#9:Z^FJbP#gG.;^M-efO^d[d<&,X3.f;J\QW&;38@U6.IAK?f
T^20C8(J/[NDN>T;2]6#D9f.FJH1b?VIB&EL]VPQCPRZGXfM8YUKTFdaY0<b>=[g
)_0-[dQBZH2=7-5-DYe[JL5]P,/M><3^].cNS6)bJVH<=5;U/KG.;H,2_U;U&,Z0
F5^;+U@g<bTT0c5X)9Z2_B9#e)HgW&4,1eDB(-G[5,OHA,,a)#L@6+<<><8+,F?G
JUQKO1aaf3N&6^W&]\,d7Ie=XF9+L=.,LE8cSY8[FUJO8XR/)UHLJ(NQ.Lc2N@6H
G+FEGKe[,=G<gC4W?E2,>X?MK<2]aRI]c/F()g6\?N#2Q-G]c,H3UbIR+6Ve3U\P
WVR:W&,>Q\dLM0,6.5=^eE3\)VPWF+WQS>4,OQ,Pd80+a#J;3BbQ)?X_4Z<H<X:J
2_.UScP:X(??T1N&0.]HE26bf0K&1HAb+I+7d9bO6WKOEH5+:G0ORca,H[./GI-1
J/>Qd@cS[^cY2V2ZOf&EV)#U6<d1Ae4<J7;Tb8F0?JaM9>W,)8KMR5WX8CMZeVg?
6)&WcXKZPSD294/3>gF@GL=ZDMF.\&R454&d#]LO]WW-fGb5J,\8aVO]5L4B/7V?
8g7N0MdL.:&Lf\f<^d[_,SZTP+M84:RM&@cXP(+X6?6Q>LCG_-+fF4c7A4YT6/dR
,ETb+944->ea1\_dH(\\OYe:b:W&IW.LZ=BC82&:PYV0ABM3FLVK)cCLF+<I\dNE
D37EOA84/C(5NWP:g2YC-=(A[fN\#FeV0]>1/5_;XV&SDc&PU(W3Y:WGL?K]]SV9
(A-eUBZ<e2-?UEX/>.24EAMeDKaGIH/UDC_/;[L?91XcEMbA1-3F#091.AD4KBVT
AWcWWS/_13L?K\-c(T],>WJ.N.8:aU3D5D:]PTOD6M?=MSE&JBKg@bXE^HJOf548
RE2]R8DXOVZFa71U[4BZU/2&-KCeWB&JVCGW#12R3BN1F4V/M+Df?dSQU^1GbI,-
JBV/e_3O#/NOKM[J:M+^N:.L9c[(WBf=Wd_/B@B22959&a)f](#K@.Y=1UMWQO#X
->RDKNOgaDN+^=,.a7A7+f0MBT^++Bd6[USQ2D0R0<&7-&=3<P@PaG>D?</?]3&S
G\?P(NE00Ge5g\^1C<9cY\HXb+gf6IZ/g_&gb@.>R@JB7_NaM1/Ce3cYP#&GD79C
9cffc&XUWfQ:2X?7[=fOL4>V.(;+?E4IZaL349,&+5]e2Ua1AO_R(@.T@ATbHRdY
1Oc2>]^_T0WP6TXWJKG913^HILTH9SY0SN6R:?)gP_J;N42@2Q0CTZB1ZI>=+e-/
.+XXS=<<IegY=@XB5?G+7J[>HRe[gLJa#M_QU=Gae\XUYSI0O;I3D,UC^\;X<>?M
7.5V7C00M&DU3dO#0C@-WBUNYVL5b#?VWG^[Z,aJVddA.L#HVVV8d6KUS6]e<U@=
I(Wa?EA1_c8AZZW=[H:R[]M4,KX8d6XGR0M=VI@U3G7.#ZLE]cb)Va(a;^=.A]+D
Q0^@f]I\L]fY,YB9aeRM4=DU4=cbCAG2TFbWC)fRPGZ<1D(3KRL-#)#QcS4TB+NU
L^I]/dK6K8(Q#A#&CHXeDOPM6aYZ1TP>D^4Y\W:_Pg1FF7U;5;<&\]@.Ub[Y3HK=
E<aHLVLc.9@XTQ.c?-VKCQWcPYMI2cS&f7T[[?fYQN_-P28WVSR+KH@>bYP#KfdN
A-X4WbJ@-f.,W=,1/6IRW_]Q\/bRCXbI6YNZ+3]DUUX,41WeSBLDDDE-SZ#>/[/M
4gK9FadSI53SLbOK8Z6b24:#FEQD1AM+))@/CPU<3Le5b;L;OdT>Z<A3?REE9MSO
[LHD9URJYE+KOg+5+0D+5B)\b8(aWc<+/VPKB)R2F4<3SH@;QEX;;fAGBA+5[:cC
4#]<KD(f6+_c3YA6BQ+\3FM=/-YH+G9L8-+ZE=&MK7BYWBLWF2d>^Y+;-Z7CO=Gb
_N[6SU2QN,15F[DH<Ug5g2/gQ]A^H^+@0>>RS18L#d/ZH=#<-(?R9EaeaP<=_()E
JY15\JOgTbG>PW3CQ-68IE.JId8cHD/PgOXJ[_B3#5PL[M:++3B4E#6J-88#J)f6
0g:<.@4P?Y?ac(J\&+JWS=0<:9AA\FZ1;Y:W0C;H=^1c><J>0BZD+G<0-M&N0?5g
A(?U\7#(]FUJc98G-__\Sg+;D=DeI\A(,@?(Wg^L,H#7be&;G=].:C>[7;SK80M3
1V+94:>62Z&,KE>aPU(N<8e/6FKOKENI4)<K(?HA:-.+O2c9B72YT-BNWYJL;2P?
(:\.6EPOEB?MS)1:[=))9A8/eD=9)W71D1]fE+)E7)WJ^..=R4P<T5,Bb)&760.4
B\)R[YH\371+[8<,1GR#A<DgD265D?Y1K^/Tf:Lf0=gH[<0=T3)HW[<ZDP+]AF;K
#Z(C_9<_4F+ccF;1;1M93>Rf=HJcgd\&]?6b,IPeCPHI[VOB/:G_f_O,)J4WM_UG
A=)[ZbDb_abB2R&b5/=&O6[J.;T,+^F1g(a64dW(>I.\@L,,:7R)e2L\\YGd[b)M
QTZ[:g4[ff8-#F#S;f?]AP13A<Rec?=NcV6PN;g:<&B)>C&T3.2VaTece,1H^e2(
GNa891E-Wc^5OR53bBJH27+;E2/>?TOOcEA\EU<>ZZdFEeX;2==P_[?f9(](J=\.
X-0a12a0<b3\JI#PH4Nf+a7ACD?E#,PBCEcV)g@G&6AZZSC3UR6G^WEQX0d,T)bI
)+E+5aM&6;N2[=bZ+CXgV,(DNC5()HH@VF<a1OA.SaC597D&#&eZQL)\TEJH]K?L
3&)=1YZD58TVOKc+^CG1WfWY_.d+BdSJ<G5A-E8Z\@U_7(VbVK&9d9a;>9GSNC/J
]Z+gJ[](?GecfdaTZY9QbbCHDXgf7K,8P+\DZ;PVZ4.DK4FH@7?NHeUQa9Kg?6@;
W]UW)49<ZOJVFb0\5W1Y8.A5@KIf)-^d^fbg.S9QI]HJ&Q=Ne?c];d-bCQF?F.&]
B\dL[KB;b2/gK&Y2SS1_>0[4XB4DBR61NT^^A]VNF=4UW(&cfZB@E&4^TN+;JDIT
ggT,_-54?27_V_6OQK8MV#2V-;U4U-)gYIKWbS79E+/NEa(<]BK7E;Rb=:#MR3Xg
G?9G>;G\ZYDCU^50.[D#<B[8YZf/4,N=9+AV:]=E:0IaRZI.aGag,7G#-QdgQ18B
,Z.YHdXI2G&c>>],ZPL[dY2U@&e<0g;I+S=-a2]4[YR=F6ZZ9Yd66_+[;F#^F&/E
<(_4&SX,4/X(5;<R(8^PIeVc27M+4Rd3YOCfa-[8VdaRYC8[TEE8KH8&BKMW)ARC
U(QF\JUZ<7@9M)g>N1c>dCEM/:d<-?I023bV&V_3Y(#AYK.2.#A(&A&CN4P+V<R/
9a-JZCeG^+WM++g6e/1gQdK40XdJRTdS?,f[TI+/&86T^D]6@)77A8_IeCCb#<?]
X;/J@]gASV/UT&R=2a@0]CK43+PJP):4,>=_)SeT9f^@?[cN8;>c:7bID<T/15bf
6#MF06[GJH+M,;4fK,WLB0)[A=0X\HZYT?K>I&VT4__ZH^LZg?:G<>MS?Q_f6f1\
N<-P)caXZ7:+S+AE(MP=;4C-[(2),/<d4I&\c3K/(bPD_8I+H95_g/7gJ6W6A9EQ
W];:e<a<TN,.W;.N>W)A7EOA>?R-M(N8UC7]FONCf>6\P5C9D=Ed2L5J?M+93[AX
R\eO5@1cR>P@F?+6eXNFAR=^?WGgF,g+M@a]:ACHC6e?2=d=,fb0..bMU]MW1C7V
/9;1NJ8)\>EL2FfE]UI]USbP:4a\+,Y\aC\EaO+:?0XPEb3W7)Z(LV-)QJ#S[IMc
K5YK;WC9>PDdN[8gA@KOIA?-dBX2P;U1,3JR>>.;1W^B_=(ZQ8XL,60OH8;,L#4c
])X62I8-?2GA^E8d[&AL;eQb&.3(80=^SaUJ1e_3<F.;XXIR8?Z0ZFOS2bKbM]T-
c(6faA-S[[H?J(T6_<T<)0<3EBVbdSI/ZGLG/ET-eX</I&_>+A:_8OXR@1I_D^#\
(f5V9-VdYO6cMdKZ;,U(B;R-E)8ZCY5<=+>ZbfXN.gVLICL00#Ba;-&:Y/)g6@a(
^>L<V>f0K(WURQ^PH0OZS4b\HQ2(6RN]CV?)a-JQBM<WG-X[6ZEeJ@4H=R];N7N9
E/5&R#[6bTa+P+)g56CEc/;6-GZ3F;O&-YRI<g+G]Ya8LNPD/PIe.XggQ.G#6.D6
F9?T=&@8,02P\@CKXJO[_6H1@P>;7.4Z&R2?7Y17HcHAMX2]\:Vb9_MCJd\Nf[(>
N<=BcA1]=HBHX>ZA3ag:d.PH:bY78\a8TV:LHZ7.W7/Pa^G^cX)-EYD#LIAW=3/T
UVaQ/T8OUgV[VE_aRgX#Hg;:?0>#J0,b.I<]L)<f9<ef_Y:7VfLd:f)>]N5\V]GM
-[Qe5#9ZDP#UV85aYA8ca+FXGB4.O_4X9.6-QF0Fe?E=;K<Q[U2Fe#SIR^2X(28W
F\b(c[Gf]OcVQ0CYa.GA@EH8TX(:+@C?d6Y>#/c:,H8N2;OXUKI6e.LcY]Pa=^?9
?)Za_9K8gNPI<N\A7B0D];3EFg5_e22-GLAIKS2S0&Y9:O?=W;7,Q\GVEGTga)Ib
W>.I:9UW1CBdP9@J5aGL3IE/=NZT(I1ZKb1CQP&CgYaf-E#)BI>Tf_KS?c9+A?5>
V/;>6I.98E&Nc5d?P5/KZS)1/X2J_U;Yd>O<aSY]?Mc;;-4_8<?VNe03<g_-IGe9
]aJ\4O;LMRUe(#,@D)MbQ(&+F-dTe1<?4Bg/B.D3HgJ),eE,;5:f#16MR<b<(Odb
(HCL1YgS73b^NB9HXdG&2CH28aa1A63Q(I5PUX&J[212=Og:1&J,?CTOV@TB91)g
0JPbHWf8cZT4E\:#W].@M;PgQ;Z[H+3F3]8<2M9<-eZ6<>J7@?PHSUDP2CIC:I98
&\A,0>(8QQWJLY^UdC:(;])]I(g\#Q/^CdV^WUF0#KKPJ_F/951S<2M^dD98<G<:
=@E5bCf,249E\e<DTMScPS6eP8LZK0C=0f.PO:f1>J&?R@a[X5N9-R1^W0eE:P.8
)\VEX[>7,D=#E<.9&50&9T;<Pe]P6]B2:K[-^[FB3dBGDS]]g9MRDQJb-4^_?EW#
W5?6Kb#62aQRd_?_5A.QHQ]J,T5TE+BN4B(7E>Zb\93YFe.I4XX0H@Xa#+<b+KO.
]IgNAB^3?\3Z[d;XHA;]^C76(?>Dg^Z5WKJ236^NZM0HOJVCE-dCdD_3UIV6R81P
>d[M#>\CD>4>?)We:=>+M\4bF=fQf98PQQIKA9XUE,1EPZ,+1?VK8NaI3\6=_XDG
4=YCa2]D_P)^LB7Y=(W;5V_d_R(CE[\#E(SWPU715Yf8LLXdKK2<Tb7;32R@6JeW
)?^eg;E#8:eJJKL(F[P6DaFM^?PdTITcJ6-eN2_b]RU(31e2IJW<2PK<EK0Rg#(S
)KW.Y448C)\;&N)N#M?;:W5+gFL(B+LZVe1^:<aPKM.2,BOV4.CIE:Re?O.42aD<
VI0W264UB.^I89Mg?FRHN[8g7;Q\/]_)5-1a@<cB;&d@LNN62+6L:Z:;B-ZXOA9H
E)\9U@CU+J?IM3Y3D]O7IB>7P@P4Z395UH9U(Z4,CgU1fU?>XZeB\QOS1BC/3OLH
RQCeB7XJYe4&77\^(U)>#Qf>[RfgJK?3#]R=gJ8^Oe:#Sf;QeR:U&DCOQ#,T9bg?
g-:3ORC3#+,)WRWY^Jc6&CWaBQ/=bQNURRRIX>D)2=KN=fM\/-CKd76]YOTE(/&_
O+V4VX9B)M_1ROD3](]L?5[(6M5G^T#@0GB/fW)K<[UYfNB8PWB(TAQ[(S>-<YMe
S2Vg5K[GM;9G:>&C7[N1Fa6<;:+N?E#/0@GHV#\\V0):-3R\.a-[T046DSOGY5)7
B3?X(ebL+=QP@Ka1#Q8+_bcdX1@NCEMDf<_-T;8/_EQ:O@&(AbZdg6&QUGQDJ\NH
DGS#a,/32JP88gcLQDGD1BVTP4]g)b:Yc[5Ef14RFF/ZOd#d7HKO?Z\fE#Y2>U>Z
&)A7KZX&JDKZYcE9Kf@_W]DOB?b.(8#b@.=Z^UT=7UJ@HY#(\<B1SSS?a>bQBQL^
;.V9MLVYe9<-6[YFeaC;+LK-WP-?C^Q,[bI;Q;9<IW@9I(6&:E@6dU,2>41f5(Sg
3IIP=<:V9Mc_(X]2242PdD>Lg#4;;/QW,Y7(JIO6>;Vb[Sd<4:<5FR1=.^I0P[KX
LYAGVV1K=[.1101ed/TP,LECO>+.E>SS1L1eUgQ]8bN#NDI#S>HI&,C492=D#Z,[
e7eGZ1[,;4L42GMS14Y/KUX^,f4Pa<PMfGYI4=9+f@=RcSO39A8Z/_<\Rbb&J2g:
,0^6Z3./UTTQ#FVERUD.1fQ\7g7]8g3:R?>aT;F\(d_g0a)Dd7\9[7X6EGY<WV\0
Sf.N>=<ZIH2K1LQ8(C:8T?EDY0N,[(A@\A#dG++aO.#(X@7[92g59R;O(.\;Ya>Q
X6/8B)8.B)G-E7HH(#4HIVI^2_cc#\aOY@2>4/TDH@@R<#=Rd]+B2>a4.TDa7Ha1
)LBAG;B&0BF_EGL,=c@V069YJ1P<=#9R\=Nc^.#aV4A-_1@<A+,_>R2L2Uc0(@^e
O5/:EE]&JKIPV2+P9;Ge\Y8aX\g[PR<=^>T_J>-#)PAHeG@=?RHFXQ]4:121EG2a
,6]2EWJNb80<I-29g:^H,_HeM\TGd3eY8dg^9K5S/^J9,:d(Y;?#6;F#NLEV/#f-
2R7-.D#QI=eIS/EB+\PD+QM\6OU,^gNcfJKAMb2S\>_Q48N//fJ?\/+&[O(UT&a#
(?:(<g4b+#G9@O^.\b8)VWQe9GE-Vb.>M/<(NMD3K[0\BZVV:<\LU_)&/_VM30_U
:@&.4U3&3M]f8SM+RQU4,#2N+.b)[P<(5DI[SFV<g#YD>S<#UZWO#:YRJEA7<)SI
gbgGGC@^#aYD.dI)6JcXdf//VV<:\NWa=69/RVH8X[_:baN\#S+28L6A20ZYZ6_D
fF24UJ>,b85=O@]2^1JWf_J@QT1/JO-+6ANe9FR\a=^8H&cIdVGC16^13d74&L3U
?A,1fW(M01R<c^D3T8>dQIg\>ACHLeH_63\9e3Yc3OP(<EIMNdU908@3Lf?B[fR-
&+K2Y^JOWHN-F3CfNUPC;=+f+&-1cUBGRW-W&P.57./[>XYe,IL\K<:-bP,K77f/
]3HfZG1Qg3J_8X<.V[d/5b9&IgE@ANC-OW@\Q:eK(Q=Xf6Ne1G5If1;T>dQ/G3/e
.]:2]a_L/QOY[L,ZJcYd2;)_VbOENB[^3ea1DH1W)OMMMZ9Wb;U2>S@+6EUT6dd#
Z:[:^[><KIfW#fgeNHH[ZYZNb/G414d3G+a1-3U,VQ[[f97eCV)7#I(8P/DWY.KS
NXWINbbGS]g5=7>_c>gb@Q@;69@:VY@T&7e9,UIVO61F8.)1.T=UH[U<b8NJeC_E
]+eAf:L9&4;S];SQ&H?(#g;:M<-25=\&8-g:+bI&7#@/f<XM]:?O5-_e(6_\,.2W
[>T=OG=5eX?b8GL(.a8U^\Y5GT^&.77Z761VRVdDKG+O09?G/9DHNWSLD1g),X<G
4f75KT\3b51?:,R033Y@e&500g87c\PWUAfKc7_6;0SEYM=ee3@<BUA7/GSdK[SH
#2WT+@<Me[K):^2VRKNLFPS5b3WEcL95ASU\-OQV,BaH3+8WSVb4J:gOZ7/TX=.]
[U\:;[[WYbKAb)MEZ^M+]0JT:gc[b7#EcSO)[BO.;S_A^7S)d:;@^Y3RC@[(LCV]
G<)1dCZ.T>J9Ed)_?.#dNR.YWY+CJ>.AM_G[&O,+T#@Q+YOD0=H6#-DX^RER+]e_
E<-TY<QP?b0gY9#TP:T5G[d73-3C5a(O@8&g/ee]5=X=]La&?;FZDb15SZP,bFY;
I:YWGb1?a>Y?D:T>6S<=24?#QEfX39XSWDAAgNcV=X&Q#687fL6cdbLGg3Sa?05I
02+cCBN-JVc57^F8EgK/E/[\NY@;]WQc?Kc[BI/6d94?X4GDM4f8O4eS2N32EP#;
8J<e0\<MU)9Z7aUc8#@SU&F_5V-&P=HVL>L96CbP&1/Yb?=FFXM<][e&U]?c<KW&
L_6Z];?/,B#9>#1HZSX&a-7P&aT20PQ\gPZ,fZf1f=6\M6b=_#1#+_D/MWP5f;Jc
bS&EOJ,;cJJ&KGGZHJL:9K5^2P#[:Z5\-P1K,AMTEUdfIeJ3U1SaLWJ[VdC&Sf(N
aO/>375I6IZBe>4X>-ZM.,HXCSgYZ5I+GD,U&CS+>^)dH8Q_M?(XTX&)&9>R?F3<
b;f+([+GB>.V)O\GB1C4N,/CPE?6:P,)8NQGEEX>47[I)1[@>&3aKP+_Sc39-UZ0
.AH?KYa[X@B#U_0Hd[a]VH+R@=?2FVVc/XYb8=g@.TY@DeYAT):24Af74cO8GYRE
D0EE^MDJ&P-[D;LSZS30WbMOEF^L=@<]U_/02ET>c4C9gSGPQG);OX6?UDJG>#Me
]X=I)9MV][ZVQCI:6gEN^C/\X^/Y.R;RY&;8;b\;74.NN_D6-X_ZV#f4JCb-FS5A
QY<Y]4:8CAe)@C25Oe6eB#.B8bBCR6=>e]5EWQ]>K(]D@YQ6L8/&N44dcN(\&[H>
6Q-R<#7T>E@^D&\bQ0gC6bE,WT<a/KE2UC/@5Je^)TgI+_AP(ce[BRJTd+I^<Z_M
RP5NH8X:2@bOF9HX)1b^SJFb)\T5I4D1U5M/gC5&(A)R:=7RHeQ8/GW:,-2.[@L2
<<Z\^T9M4MLPb9V^U1?J6Y:B7I\(1]RAX_A5LR)<gR]KcV3C-#W1J9gJa)NDL2ZV
KAAf+5bP+_Q\I1S6E&0c/.-D^MG4(<SE<cUXX];K3IW(6Fe7<F<>,:b#SU^RA_Te
MdQ(I0_N7]?MQHF;H)_0eJS&GLIZfbFYgd:=@]#3PZ@WH[JOVUf2TK:B(T+<4AaK
70HL@MP7X(-]3Q]M_b:59WMB:P^9[NbWA1PBNW)P]P3aK_SJTCD8?))+gYMf]2B>
?+\ab&9Q-IB+;D>_42CNK:8/I8=,b@X^+LZ6@H3;0aTKf[31^@N2[YTV)g^d_Ee-
bTbLS9+\Nb>eL#a=U-N3:D?UUcO1L8WX/(\LRG8MX>UNHeYYe2FUa]g/S&O0KRJ8
VFB)FMC@,+/BN;.<7)KWY6K=1NR4c/bW0V^(K>ce8e)QBZ]KKYYM(GVS8G8Rb9M6
90LV#@H9>B#=<MeFKdV>_#bQUT,2\9]b;d0UA^(6#+a.3\0Q(]A&66LgK]U-TNW:
/8:S03V6Yb(CU]@F(.?/7J8UeeR#]O&/d;-<_K?6cQLeZ3gAY.+;C7>1[B9Na5M/
d23I/#?S6-?)&0c)b:TIY,Fb)SB/^[=P1ZW8UEcBAQ.>4b9[8?T-X<X.-#OZDN7=
2dQd\K2VP0,GFT70IE1,VMf7\e=7:0MaPcMY4+&MK9aN&gdd6\YDNA95E1,,BcZd
0e9LU<CaK^>_?3ETU7LNB#e#[3-9=1#V4MZYIYd@9NKR.B=)b:Z4PdBY/R\/?aI[
[ARV48,-ga]NgR,fRg;-YZ(Z?6>Af.e_#66N+0:WP,cV>QZU@gDX9F.d_?\Sg>=L
+Z@C?N3?edXTXR+BJc+2JD=OV3PZ_G=2<)aH:UCe_YOfQRZ3C2J1EB:PWEX&abd2
/7ZJb4PL_&V3O,B/Q-gg0U-CO)-C.JWB=>PT[BE(>bW6Y:[TP)/bFaR;c>Wc:37/
+39Vf]J+a5?]@S_8JK3SL-I@A54L_[\8N]XX./^\PH<&7[C1(gYMW(KHP_AD2dR;
Z.6V&MO>DCbX^0gNUN\T[?A=JH2?F)fS=KXE><7Me=F(0PE#6a>Z,SB[92P\;d<5
J)>=/LM,(H#NY;3N=<S(_@+(PGK>?dQT+FC^;P&:P_EAe5,JD/,ZFX@&CggHY4Ae
D]M4&V5,Q_3^f.CJZBf\=#CJNJ2Df(U+F+(Y+6R_gUdN440gB-\3U.J_,dUgFZ&9
\SMA+W:ffQZL_A6@>a8EHYc7d6.YUJ/Yf8OW3=S+c+8,T?QV>8W#KeVb4BB7Qc#^
L@49fGHO.Uc.[?^BN..I\d?f7^K7bWA4AIeEO:LN1U8]^A\_FCSG-F/?N6b:.5d1
A(NKN<1b.P1KK-\E0D9)GJg(EL-f-a5&7_BgTY\aCI,@PBWdE8K5K^Nc;d#I:+LW
HKAGF23L\K)\<)7AH]&IKf@EP?:La4Ag\.8eKDVQ2M/XAdGZOUeT&/b_fdP_.QOF
,TWB4IJ;UG@.HbNc2Ag,9_BB)7),X6ZbDM=<1@)4W+-5a2IECdXC4@_D;.,/cH/@
a_\C8-G:Vf^H[&e#2eO/9M(9d,.><(7K-OKJT]@WF(SJ&>Z@@Y&+VAP62?72K?1c
f3?MGZYY8T==]fYNC=@IeQH;X,a(N7S_OQJ3OMNZJ8NVDSX;,?A=YV=F,C]Zd\BI
/JDIEL;&gR5<N5XQQ6PL,:<=Z?-b<Ha5U2LI\K2N>M)f@C2YE:FPD?[<.TTS6ZMb
<G@/\I_G32AZ8Oe?XagHV1YS@#c0VCeK#ERLP1bGDIW9E@L&9SOM._:Da@9?AeA6
#PZ#L7G&_FPcVAE4O#]FK],R4a30VbOb@aXSc2-Q_6\<bC=)VH8OKJU>>BV>\#V&
7L6&6+^BLX(QD&J.1Q?5,/XQ.@\#cG8-[H0B/19&b?/IU41Z8./0=fS6N/DcR&+3
e;@8E@U.),+a[L@1\Fg2V<JNdeSI<G.d2)K1B>]a<C]I[K>QC@UTRY<O.6QT@P\S
9V<82eQ.FA-<IA@M&H@NO^^5f@B.^DF6&Z]6=&bW:YGX=;XNI,;c5bO0KBVVc&<;
_>8<HL+fIc.Q9&37eI&TW3D.20dF#)90&#36]+SUCSI/D(VJ7,2&GB=7/R0:ZJIH
EVSg2U^0[\0X]DZHU+aS(H&cE.WE^)5-ZEPQI0J/KF[]OOC/RL:9:gEc:7aOZE6g
=0R\^VFKK1N0Z0d3=Ae8gH>2>MQZA&@Z_2H6VPRAV6g].L45CRMWYCS<bQbYG3MG
8LJL?>c:A[RSV]QbI0_6TaJO.DH-8?(0GSZPW.E^EY+:Z6V&232>7D?68eg3gSFV
0e6F\;[1M=^RQ;7B0;bR:3V\M0#ZaGV,cgU<_PAc(-2\EdZ&@1dTCGL_V,AI@/HR
dXg.A4NH/O\]<V2bF?9^3=HMYD5DEDQ3X+4^Q(M)VN-,_4+:JUXQ6BfYC>bK-Y2)
,g^YdD9Y;@IPMNV/8f9SKY,G;?Kb8gQG^:d-PMSW:UVX[K>VG?Sf3aKbYQAD\6@D
,>_LZc<.B0HZV/,e&0cV)3_bLb#5O>;:UW#95[aR&&).Cb>2))W#D8e\gLQSfb#X
S.1J.a86N#TU]5d[_397]KJSY@)KW,XF0ZAFC/:@C\0X.:5:=/f+1-;aTcT>H(SI
:@B^T<X:GM+eCN1V,\TOd2WBRIATO->GVUL1TDG#:Q>NEZX8QG]WDe9[QR&9@Tc8
67L7J1XY\T[\UUA3(DW9?\4/J&.TNX)KeFFT?a&Q+#]:5,CP@);2G^C0^Q8+bNLP
WEb-WJeDe9?+dbbW>6#Na;e.])8@a@6/bENU6,EC2J&cNE27W]U).>&IM54ceG.7
RA?1HF\/.[bS(EE=b:([M9[C-B>+L5+@OPZO[O0H49ZD0AJ-@P()IfF5<C)gNY.f
9>:?g\Wb@#3R,+-D^\9<0a)R,(aPc(60),2:I@K?6K=QcEGc>d?5@ND5a-@GbHTZ
GHI7&DTg]6,YAdWI(_BQS_\O1@KN&GIR0VUaG[3RUda7)a-N-fe1Me,f1.E3\aVM
KMa#LGgfP52J#8J(&(IY/6Ne:69@HQL4?^IX6LZ>LgD(I8FR:R85LZG[@fF26>T#
7H:-SET=e]5WS2DN.=A(-/Z<6OVG&_K+AR/=2=0Bcad#d_Na1S5[O?Y6b19,6F>=
)gI>409/F@5Kc/ga,@:BUc)QVRYA0G4e?fad?@Z8D#71Y?GdP45VA8S9RVEb_.[1
>XD7LKX@eTNX=CUS]\.Z7ZF^X<D[3BBD]1bZFcfBd0JL\=];+RI\ge442L+(LS4Y
-&=I>B>?,T\?:0#4CO=^R9#65X8[bW_-.Tg?)4_+JQQSQ>_;=_IJ7@TAK(DBQU5I
DBWbXB?CHA3;LC+MR[VLEegQ)99J)I7,bA?Y[efMQB613cQ?:KU7<IN]KaY/9<)X
I).9bC6N1-;K2eCEX9S<P7H4+H>YaJ4#H](G81RI)>8:4-cMTCHC&Z;0X=(7;?6I
PJK>.^N7<gWWWG><MJ15\eK)]dF#G_=L_7fRUT85=R9cJF[2Pg1ZNX5d/VJ<b3.c
-#^bI<fKJOR42NgHReZXgP-eYQZBN1Y#C5S5+[^Q3>+>dI6^(0f6c.0CV^TN]:,[
5RPZ^U1V3-P#G6>]>C<OLBSHNA48]+QRVa;+)]UHH[PS\2[;+=baC3F,cT-(A,]c
8<5Qa^D=D>gE3EBgANN]+fZ&(V.+J[e3a>DP3d57GKBf6c7/?\_K1L]R_F[2AfR3
S4;8TE7+9Md/?LGeVeJFPTI+PbbA7ST>SUWMQZ#c-JL9:J2R6C;/;K3;,F6KaYg/
7;R8g_N#W)DAB0Gae-:C8a5_EUB<O[Y5NA@1@,3JQC)8Vc2KM00?UN1^Sb&8&YfZ
AKSTED[P^-]/6L/UTg?1-Y[OW^ATL@8TDP)aZ7B+D@O9]M<@R;&]eEL05TKb4,T[
0f2aAa8]XWg6c+2S0^\6TR1NDV\#NU6-6_&-_IgV>5^DVd3)93^_K_:HDGE)56Hg
H#ae>Dd]c_<LW>VQ4&8@-\&gP0SV69+KDM+(XK7OODHLTNXNCVVS6LCCbX(-G,^U
^1<gJQS[a8W&c^/0.XfRGT2^>6K(FTB6/R\ELYKEbSeS.,_IB>_<_FV[5=a.]@[)
[R.VPMA?F\B_.B\:[Wb-\/T\2I(L-Z;^cS_M,/UBNJI&9S&E2TeIU,]-^F7Qc]RG
BgG0@IS>QPaQ]a+JG4F,#BaD0Oc#A<2GJa6E^?VTFe&4^H.\:+H.1Zbe1R0>?YCZ
YP_^;2YC,bYW7NI.@@9d3?-1eUJS4_\a<A4>&29.6@+8-AO33-80aRUMDVJM9_HD
Z\A]6I>-W9JTRcS6A5?I2ZPV6L;4NJXc&-9E8fe<V0fOI?MG=a)6fbR)=KD-WBfA
:V6L1K[2:>f70_=/YZZd68=K)[#,.M9.-AA]]=HBPH3Y0eSQJ/JJT,Ce7(VU<&^T
81R.E2GWQ=3DNe7ET0?+M3&H(bT;5a>a323e[0/MWa\7YWa@_.;SG]8QeQ<f&ZeK
H>_ILG-+XdR:(+a+G[,H+1\[6CZ78[N2CQYAc,L/64Yd\XKPEPFL3TU@aS:EXFT/
7<Y&.8RJeG,\&f^Q_<GHf7ZaUGG#Z.[;7JeZX;6<4JPg_L:9,SI:=L_2DGBC-NCd
R&,g\/B.)\HUQDG;KKD5Z(+[1eCL0N.,=;+BfM?,9[[64g8G)IJHGFIF6R:N[P=O
&?Ze4O2Z_:[WQ-<+4NB(L-4[JA9b5VQ.8=]CacBH9NZ&aeI1C@U)M-cNJ62XREYN
JNBNMU6[:JRV7U0+]?767WXdG6^JAgOGeTB7=UX2FSF/KAcRDYJ-Q3W9#8J,(53,
QaR,S@LZeN;C_+=C6WBN,BH-W-+I,P8V@NHUPSLRJZO\[I[\05?A#b<XfHf[/=#Z
>3cFDG?.IB+cLI7V^IU7A=:(J1@V@?(WUB^?@YPHM+8f;#gP)NXQVa(RKAYL8d1?
@U(A+ff>,+)HZ&\L[@ML,4@bYGSML\3<KTfeB86#]7d?fGTLA>G&R+)1(\.g:173
D8):A)T,+.J-ITF[</-NTMY^#Of#5E/5^WI=[ARTK9g8(ZQQMT^E]6_O>QBO7g_3
J6_JgC=G2WO-QATAT9@;MN;1Ga6IVN2gbV;9K24PK<&:X=L9NL:#TJZ+)e\W[A>T
#_f3BX=15K8=_(ZWec4&7#\@Ec10#S\Lf]S;AC9ICb(7&F69PE,IAY-X-f4e:64f
[82S\51ffC/=3VBRVR.B\K_]A>Y,;Y+SNFDHcA3FLcV;M(]A:>NK,^c[a500gf]&
L\0ePRDP0UO]e-UVPeA(ATP]6+R3]=.5V+2AFf,[26T862^3g4c78a8JN90S2VN7
b=6WPAcU[ECOYP5XT2Pc)g0,6SH<<9[QX:2BWO([O8N^\23V4)4R@a\bV2U\.Rg-
fdg9YA>P<:50DPA.+B?HA?J^@4gTKV[T\E--[CG^YT+83,J.D@1eV2#42f29/dO9
N2b2-8eP,,-7@\]bOLW@<=@@5H;4M/<IOF<8]XT9991<99Q(73V==4M,9UTEc_,d
C]^7)1SS?4#9Y)R&TU/MSX<eaagQ[3JQ4eJ(0J]LB4&)JOgF<3M>3VY5,5G(Z-Q;
R,LRRbEb_<)HS\S^d5:-=Z4CO):E0HcKUUZg.0)2c5ZgR)XXc)228U8959Gd0295
eEa1Aa-Aa9B]X)Ue^FGSc:UaV85R^Nb(-@[C]@QOYHR_c1>LN^_^M/64]9ga-@Ud
7,GgMHD:M^?E\R,<R04If_^?.&U2^a2&:T8=GE=d-5JeceAO)PZJg6P+G[M?0^cG
EO(/Lc+^99YPQ-A^>XGG_D8[[U+N<dC6ML[8#ISRa+\8+4C:&2R&Qc:K^Z^LCfYg
S^B49S[]VY@dG4<^W#JV<2N2TGVGEfcZS&SYa;e;Gg<Z^I>JS,W7EJE&dc@)1INA
=32agYZ__PBM[#?P;;_f[46-J-?NF:>GXV-Y,^^]1Q[3-/]UZ)LZ)I&J?:N_SKAa
LLe\T0<&9#VUMTa?HIAG=_V2/LJ)Y+1PD)Q/PDNN@QG#5LC=G9^R]5FR1>g+WPdg
+[WV_JeU)QH&>HU^@;-JJ(L0W#B<@0QR@H45XF;PbT[0(2)>)X6-\ODBd#:bJNX=
c&:aM2?b-d/ed#Z2]JfCLN)UHAR7eIZHM\GV;<d]QS?&OOM<6UKS3^O]6./37>_J
UP<]+aGD#2c<YC;YeG&cG&+;Rfe911Og\:R&/;4?0LI1S\bc^[U_:a)&FBaaTOEg
&\c>WeC\H8CQUTf0PYDS.7@JL]N_?^2:1(&/(gfc:X8ddb8W04c38:L&4&\XY94.
<R6GCFY\6aP7ZNb7e[2TB(X-H3GA2+S^Q<#EP^&<#]FMI.4T6,;55M/_X&ASEA]f
TD_Fbc:1O[SWN.G(acb/F>dFMXT>f4G5RO<S,bddYFf8>S(HJI1@A4d8550@WNXW
dKNJK=;N<=;S#&#E71+</f4dN6:QHFW9[3QC1,T=6eW-+8B@;3bXO5^G#OAb,M,;
I3Hb+^1OOCZ[-#F8&E,)D5@C?^SZT9e[<)BZ&43UY4].72bd&3/T;^G5cO9?B#K1
=d2=3gOYN5DaNU[5N,f(d]b<D0TV,9UL&R1^2g_:&dcQ+GN+fXD70/K+I#WWCd6)
W+O.)cI@LBV3&,GK>@#CBb>.FW:Gb)LaId5:@cZXZMOa99Y2\6b6[C-ag(0D>E#Q
--=KaVTSK^dW4+>1Qg1.OLLHaVS=G+Q.SW#1G5DRbO:Z(:.1b.4BXI4b5,T>_CO<
H7-Sa7AGB.Q6MI(BC;W]HfT[##M#dg#d],U2@[Y<(8R5S+0.[&DTIe0<D.IEAPOK
eF&4+D-QGO/@[O#/NV7XIKf^A[[/V&?814K3S:8F6VI5&_+)V+_-#J#A]YCIcM1b
R8QdF/c[07=\DR,56@,[N(,-ea7/1#,\JH4;AgX3fUBXJQJ9Q2GFA<UfPO4:C9^S
[PA7\#REXa+=6d],/UCFKU3+;O=O9-d81(:=.LZMR:9>dCQ_2&U)&GT4dB=,W>LG
2=+[39g&f(CA\^7##)bTc9E[_bG8aaIXAPHMfd\Kg;C]U)aH>+<P(_RbUU&YUX2:
FVIVac,GgcacAUD/[A\89WG^BLVc.=(R/=)b,M+P6]Zb.^,?/f>7VBMTC:A.\?OI
2T_&f8aW/1E9GQGf2JLGK]J@\6bW^7HHd2a]Y)?.-;@MYZ9,GP/I+DDCdA?R<Y>:
9)+H[0(H]-Ec[-0Q<^)X)aSgc#9X>14<V:ZCJ?0/VG98=ULU,3f@&(BF9].9^fB+
LS#8:6RVV]]6UL#Rg151QRU=EE/c?TM6F29@2c^^[HAGg@7Ic&9</?Z-E2T&K275
&\c;VNe3LI#U?-WfOG=Na7-CC:S5.ae5\eOf9f:3FBcHX)<VX;f0]1_[A^P.^g@<
TCG/a<;9E.9ID<,YBQ5cE@3XWDdKDcYC;a>)abH&A&<^O#gSA>L99Z86NCgT[6TU
Z,IOK1&<I=]7HaBdEVP=9=1Z;98f8=aGKF][HE;N?eY7cX,df5I&XAAY^NSR?YGA
e;U-W#=;AG\:D]393;C2fNCZ9I1RF=&:Kg8f6#A0S:3D-/_0?&Z0IV&J5]RS3]M(
SDI456O;QHDN8-NRGQ?&:7:AEYE3d-(/e^a&HX2Pa([6bRe5^6FIF>DG+5#RF3?>
4gRI(L6N.Qa@=#dEGEeaRD[W^S1>Ya?+Wd:,e]YZ.<f4bQTR<>UZ)U:@6\.aZSV=
I=g1d22(gWCH?f(JRKSXQUdHU&9;=_NF-S6R)McRJ[L[+>FXA))Gfd(&[NO#845[
F3L8@#?He.Y1fRHP>3ML8:FUXOdQ5-4/=W25X>RML-.Z&[XKgF7e\S03Og,]DOB>
E\=5N[^QGdHX]fMD\[&9D\QG=VXK6<U8PVQ<-#@fG.@T<W2U]O[63[#2eI6;Y;>e
@OSB&_?ad#B)[B?\V+8_QV>?OYHXFM55:L:?+QTXO?#9_P5Oe]_U?c7bZYdD6IR3
=SMNS<M^IO=;2Q64abS]HO\NZa[45VA75U6]FPa;;DJT]@/80Y+&Y,&H3>^^g#bS
.4;8>U:#Od1gZGBV4#T@<Q)DTRa#9E]]VPDI6(D6fe2a[M\/B+UPDC-8GI90b=_;
0E4#4GK3/+:PD+PL48Y<+E,7.:gA/7ZX)=MK]=cfbPMg1Y=:I#WGa)Mg[)GDS^&G
LHe;59b2c5_=9RP2;UWW>TOeJ95PM]1)VB6J4=XIT([X]^5\I3gS4ggdaVPK#0EN
MC)IG7IdXd&aL]QP[4(8E&A9U=XVVR.e@-gBA6ZF_@cZ5ab8fX&1c9PM?.TM?==D
cB)FUgP[MN+#W&]3:.ecU]^1P]D7)fM.6B@^&HdTG;1D:e.6Hd3Oba\8(+--;S?f
8(A?Va4M=N+A&1,:^A>N=,42\^>Q\G&02a1W,gcJ1>[<+_S4K-,c3\V)&L8BVTgD
Z1#4WDG\^;FgSQ:MY5HFX[OC[01B/b@DX+\[/S(DD.QIC6Se<T]6#RZTaNDeN91@
>]MMbH<3gL@-<7,QCaO3J99N2LV,Ue.H/<JU/6C<ZRA:Lf1@JeIaP0;/07aG(4[,
8TFTDL2J\6#3V<_X<9fG0(QCQ>/5YR-2[R.Y/__=LN=^.eP;D8d.ESDJC^2eJ;XA
PSDd>DeA2TG@?&>J4)=Z0^ge+V2[#f(+TI21f]dFcFT(UONZ<[NXYPUB+<0e00<I
IfRWcW=.B#87+XcOMaZc^V_SM+4Q8a)F)?<0e;FJ1>=aaW)Kf[=68(U]\GZ)HDCV
Wd8:efMICFADaaPXI#bAZDCfHP8SBbX=89CWZ08JBO99b@4?QYY+GP9&5JQADE]A
?Y?6a2Xbf@HMb57F7R04LNH?6BWO@BN^2W93JY5;T.[Ab9GATV^HU@GD)-/g4+W)
5fMBbbA;V(>QEfUMRKMZZ,F=e?,52+/#Pe;bI+3YeGY3Q._ZfJ2SPIWQ]1C8GJgC
ELaJQ\=H.(J7K7+RKGDX+#;=>5N_E))VR\)10^@GO+gQ\\D51#E48B]TN/(;?7=N
Xf.[fK;F(:T1MT_B7E0bXJ-/E8&5AgML,NZXDHM+-C^5FW<UOg/N0KPV;=Y&QPAX
0f>d:&FIS3a&;U#3HISEM(2T7;17f<GCL9.H);E;Ra=0CF-[UF.aFbHeb)QJ0YO/
3^VgO3R-GB3gU)/b,=UT3HbM2dgScQ=YLQT>\BBXUc0\]bBM13Q:D8f6SWaD_6^#
9_-Na98^H[Y=HCS5F3)P:6EPA=P:U?XRJ+>&0XcgA#G(C+gL?b6>^5U/+<d1T<WS
A7)6]QOI=HC[Y:/;Nb?G3Y@B6-3#Z=c=3BWd&8P@-7,YVeRNdK9]R_AMUE)B;XX&
F:6(+?\B7[LE7bC9aI#f-,]=P/c]<DE>HGOX:O-/]UC#S<P5R0+?0P)H&Hc:1LXA
5.9)25WQFeJJ3/bNc08RRXOR;^;TYNR@F@QS.W6LJ2EO?]Dc/3LeMBcg=81:E;aX
ZSfa9;Q..526J9A<VF]]H822H;Be6]:W(dY:JJ]>V^1Q(+3[JE4+IV:#R#;(5GA,
5dbPBF4EB2?(GgdT<g=1DSBg8+EbTV\X<a=PE^AN]:40#<\RM0]7^^]R)D)&68;K
KKVLM\8H>@QK-25gGE^)2RKGeEJ;I/L\.3.g2+7[7Q4\1ZZRTPM<RJ\P7I>,_cdT
;SVVb=9TS8/#Z&<aN;eKWOTcWE\B0XJPWg]2BY.;ES11O5,=J]1>,=3&LR41#C[X
IM/4.Sb7DIZd1G<NKYSE-aP3dZ;)??cQ>\/K/OW7aOW7YA;PRD/>?dGd_TF:1_e6
/P\-93M6BU/aW:cf)X^eVe?g8E>-AASP?)@-PT9:Rca,^OA;L.M#RUJ5:@>-Da64
/N(_5J&ICP^G?e1\]6&W020Z:CD7)D@F_]F=dRKHO[OcP.aQ0X;57ZOH;UMLH</G
&^cUX4Ub7G^#4FR3IKFM<gg6?Z2IRKGM6:\,C^_BfLMc(0/W;.L7<93XUdSO9\\@
]#@I7,a0PFW_RQED1g1Od,(N7<)U5PHN]f>0,4UZ62S+[T>XD;@CIfS>>IdSZ)AD
;?a=G4Ee,#b/_HF#Y2dgHC_f:DWTX>0050KJL)AYSZ(Q^7La?S2bPf2X(J_4RR2V
L07H#,COUL5>HR90MYTX,LbfZdb8NR,#LO8H6Ud7bS3@<F9d.e[J5df.Y_3HOKK2
/dF,QKLUK=[XP6TE0^FE?e=gCI/,YF<IOQ?5/-9W,6<]g-K-.&TPL0gEe4fc?:NM
:ZBV]MU:=CC1CGPg0V[HUXI&W-W=\g6#?B;.YUH=_7:;ESXYS?IE+<Mb1NZG_@cT
_c+bT_)F91M+,bC;ZS6LI9JBbbSQ>2)0b1aO72T4dU2N7BO,[A]YLT13D-BMQF>X
VG6E[Z,^YN(QTRZG>#W)@;Zb\<1NGYHD@d<aL>f<JUf]gS\)6WS;9A<_NT^<4UI+
cEXLE^cb]b9acYSgaVEd(FLO(RX,W@M(G=(2RGEeJ?:I0a#O_S-M,;\gXLWAG>4K
CU8NWXZ3/HWW(QaE@YVKc=/2MCIM3ZNBP3:6)OK\TM@Vg?3PY^>YPW^&X\TT[a15
S:MW91^\AVP[3ADcF9KUN/[VT+KX]WR4ER9^Q[CPF4#AP4REAbCRM[RS7MS1KJeT
1E(3E-=F)5M5a/1,[ZODM48?01Y6KbHWBIZ8</:XVgYOgB3c3&I.0O92(Q/QcJ0;
VH\U><,S^U@2e/5VNa._>BL^>>U0QIXaB)<Q;DP3KGML[f7EFfMU3TMPR+P3O.dg
WFPBVA=bbKC]>AS4.8CND<1I@,d1W5[:ag9DL7EeL#.+>@2Y\G-IDg)=Y&C@R-SN
W#WHUJM(N0eBEd_>PE>N@#>S8,K)/_G4IfK-DMV&RB^G(BLN#G5fB=/?M+[2IS(&
@R5E:cM7,R4.;O9&&]1=W2NOY=2@VYM>b4J,PCL0+-&0dP((<c;HT5.gH+0TdHG[
>^+(2-D2@0G&,Z[A3TE8.=U_^XS/T]6Wf<R=bS[?e5MTN5Ya<]0g[/3KU,3T)]1H
+8Qc>MX.M6Pa4-6b7SV;=-T4LMH0c\2A&CAOJC-<YZ.7\))5R+NFR7=-/RIaR@W8
::B9+^26^L&,L6F<^[O2,9g;/C./(aV>8+-=/dVOY,ZR1K>R]H4V]YX\MeBR<G?B
d8E=VDJe3UK,=g@O<(gDd/,O/)7:<U/>(fU5Z&dVOcRSTM0PMXSCT;X\]/EB(bB_
UK:6aQ\XA#PP#Se^gLQ2c8V)G(ADWOE(RAE)HQYIc-S>Q6^WY4M6L)/-X;.7Z)EA
&:a=g^(I.^,6b<eE7SNA#+Ebf/8>Z^PS;7/@HMg\g=_gZEZdTCc.f\D1E)H,H[gI
\eeQgX3d^KDKH2a9cFd3P;S[\+>7&NdE0Q[B&DU548CM8U,BH-Gg51Z,;55BLG/-
PAWS?2,02C,/6J?V4=(SWZ):]9<E8d+)5B.Y&6?52:78C,WERB,F&;K#()VaN;.>
+V3_,N5M/QQ]?8gO+MG[-VQZ\;-:.96K5?E\],L]5,J8OW[f#5)Mf/:g4IHE+P8g
GEW]L(4QWg/+_&,PVQ=0NP]__7>/O.(4-gU#X0@7;4@E^P7=F3Nd/C9_D:c)eeYQ
&dZf1[-YI;<WL]VCV)M;EeN,3?7F0b1<]g(M00A2-2>PD[GISJ854Oe8[L8fZWZI
eH)bfUCEAdN;0(Z<dO3Q1U+(HVMg6Dd3d[@RZ^=)0\OF[+\?QGC(f)YK:d6I7=EA
L3&?@DNZN>77e]0<AN+gF)APFc(&.fS5@Pd?866a7[M+3+()Y+_XGTIQ0<;1KW/^
),fg5J3.1.B\6fYR-P5U/_\95>,79.fC4E+9G\VQ^[W;3L=S:D7@6P\9,bJ627Eg
4.d/WSEBc^d>65R<Y)g5UOdOX;N0D?#)&J@Ba6TXe[#FdJ5(/YGDG6KS.2^F@?E4
\TG&VQ]C)VOFWfI/AVEY2D6e7f/Pd0<#d1IfR#@]UTE@AK&L7N6YKg6W/+KO+P?b
&L>4H3cIU12IQGH?P)HP\G0LSB+N[-10PDXEdE;O)e@G3RGF@H+dS7>5H7\3NJ]c
(=C_HC2VTB_P&Q:.AfZcF/X;K(#S[OL.LA-:T3GI>=^f-1-QL=BU5G_WNcBN;gUA
[D&f4T?d^=)_=f8/92XLY>ETRg2XFa=:&AP&+,V^7;W&2gDE;JKc,2RA:##I0DMZ
/.YH/5^#bgXS<d+(9(dePa^X]?9+YHO@dM2E3JS38SAK]@D;G<L5.L(8&aHY^O\T
66M=8JPJ;3,PH^3dRT2T8&RRM&gCF+D-FH(2G\A88f[;8:;@D.J?6;JdIOaf_0SN
53EX=B2H\&>c[/[:K;7Kaa[UJ)>KV[T#6T?#5^aAIR\TE0\D5N>e=#M.-B7V\e>I
_g.\TGefX^fZA-T,TA51SBG8[AOI,L_=3NMB8_LG#GWVI;8/H@S0>;82\48XLKaM
<N&MG#(FMQ3?Md-UB=;SDSZX9aQ-I+,#Gf-#c<&(dXYOfE#<6M<Q+UPLM.(H5;+R
.g/9D-@DR.)SIF,?I4eS>C\TbTZRGgA)8J3]^aFa,9\5B,c8D)<MXVD:Dg/b</S^
\IEEH)TFfI)#3D9ZFQ=:>--7@2<UdU8F#-:/FIZB;+c<B#a;KHLF3Q4V7TUHG=_4
Je2/&g\9SGO1WER>[J8ZDA=Z6@CCOI+-^DVE_B]+LfO2(1f8f#E9H4/V[(>?fK+6
,K5K3H/XR>1&HW4\72[17f;SC5M0Pa-a6)EO0[J8--6G73W8D3\E3\+<e>_Lcdgf
A9O_(+3dAM8B1AS,@(]_0(1,;5G.K-C:/2^-Yd,_9<-BR-aLYFV&^ZKH6,=&-fcH
g.CHfZU8+2LN.=#R^8e-XOEU#<#\/=B^+>1a^A,S;F6ZFO.B&],FHY#>:NOTN9JS
UCLZB#60V5-K94LDa:(#9Y<_b\?gTcYN0>:0cb4Y]?G5L@A#,6?F)_cTaE&^JeK]
_N=BZTNKHC2dIZR-f(+I:d8(@0&[f/]C/+GXe:DAREN6X83N,>PSHf[9?0=;E7VY
AY?=@+^9IK;.8/]Z<=S6a4c8aDfb:@6_.WF/X7U8.9=d2\:8aE;Y8J]LLF+P:UGb
PTg06=@7F^UX^]L>ZSQF;5,1f)A),Z0;>NI+ZVHF<0_358IOfLfYa@<dP#)3Q=,U
<.Ud[>R9QK670+LRL>LJ-#KI.gVa8T=4^QU>8=XR;NY-WI9e@L/4d-@-[aK=B=UC
.Tb;+CZ0XeFY9c[U)_-:0VdCN<VW+>3JM0:Aa(?OKa8ARD+V93S)^IMb8\;7X\JE
?FIOHC7AMb(g14+Q-C?J_c1=VF2LY\K4^PbW.C)[NIR^.,(GZPZ>?294E3)8eP3X
,9B&V\Mb>)KON<@87<^6<Sf(:+a-R^(QR[1_J\[7Re/Yd1:b8dZQ4#W2;,>,=MWD
W#5DIHGA)NXd65G7-#(+9Q(E?@/[CID/4)IM=MJ2-MUXXL>,Qb<RV0/fEKTcD#[;
cf[37b\Z5JC@^YV9EfaF8YY:3#EM&caPL(D?f^OcUWSO1N(2Yaa;,<6TfMP_-bUJ
[e4(=9<:bSfNQbg[#MQ/[JZG;/fEM.)5PUH?/-dIVEf>ecaR[E4MZWX7e^=;F6H1
O?C8ZH;43LP?ZcU95;POP&D,6W]83[e,&MaG@A(;[0^)PMYR/O@&ZFFfZ)S09?5g
d(Y)d:/9O2@XOZ,PNWX.&^MA2F952<0eLM8<DBM&ddN^>2)^0b[0W479@]ORR[=Q
.AV==M5?4aQXXY&\Z=8eg-0c9W)MV=&gJe&RWa;&J,I5G2/34;X.6AAAIC_NU-(2
39<=J_)=KH^B6MNBHH[USaECH<SNQ,T0:=4da;BQT3BW@4&LAgbYEX:.0)4#)4I6
<D2VJNBbI&9CZD[XUXMT<H0N)84ND<@#O@6e7A/8U5:O[cGAU];6Lg:JVIf<EVLD
/1/cJ2+99XaOda6?]/V<c]WJB?K^O;+\b2OK2ZB2c3P[SS[+P3C?KMM1+A38\U_^
6PMDZ>[+,1GW,CN@3M-f+&,,gGR@D.FQc0[[LRX)1D)HY<8RcaM/P/>R4@3>XJ)M
#TO-ef_WU>BS&NXbP#:8575_U9B8dI,C8-WV?3LI5#B6&fT+\2KVSROAFTP141g0
.PDcV0L?S/;#^+S&X1S4CZ1DV62SMUN\\]/1ea(a13T\#<EeHe.]Q/K<J2@K)QPM
>T.Z#2KMOT_39FO)\TX@3QgM=c2RT6(C0B)3D@@)W=X.:JG__F8Tbf8J^=+3]T9R
71G_,UK;&0eP79#fJ#4^CFQ9Od<)KAB+4EGRVRJ-)FVTJV>]QWV6DUABC?>F;]-M
b@B1>aKB,Gb\4):N]5\5)IH#O@dFG2ZMZ]7;.g6+C/R=YMcY,=0.\@JYUXTZa#1]
>VN153F:^6Da1I_ZKVAdMK/a@3XD+4L5W219>3d\#V#1DU\UA_0CN>&K=8Q3<K+6
@JGZLB[@-6gV?fXZe(4>)@)AGe1J.7<fO:C+Y52>,/+D1HKT4FV(W9^^EeC[(f7/
(]2IA2MRY\bK:>,9&d).9?SGT\fZ\+Q4cUKO0bYc_CO>c5RQ9:d+<Z&US6KYM;?c
Wa&.@WA1M)PN[8NE7[,ZQ2^Ac-F\JU,C(78@IQ6TOL/+dMSNOA4/Kf\GGL:HgD@T
/-UGe7:dJTFSRbPAO)/@?CdG]>.+QY]ZVUR2<e2#B&DUQK>CZC326S2N#U6WRd#,
I#D?H.WN#JXE;gg>N^1/:1-&<;,1/\6@,7f:G(11-caSTf1:Pc1VBIA]4A;L6=0K
b6bbYPC^4\7fZRf8g>4JJ:/e?7+-ZG8ZC#IB1<)5C?\,P1XHCAaH59TF[:@3[9@Q
?f9&F8H&aE5?1;e>A9OPGNAWU424AAU]5g+I?#4Q4JFG-XdLR_T\5O-.Ag3=^+de
N4J^-a[SbZICa83B:6(>Pa2)dE,OBR&/gI#cYL\X,,4:CbYCG81]3PKOKD1QY&#^
)YL5SQ:S48QXBgXOHf7<SQY<:_K3:1^X#)NX1aF=GbF^5Q,H>R(E?>7CTRHEZ4PA
QGb?5SW8]I#UdL3NZRHBTMC602[:O>d\HB(=eDEKETLaR0AH:1D:^,U\/X@L&[;0
Tb3@3Cd,(O[\DAS:BEIX+[B@(Se4GSU4\/9Q+H272dR.Q3>&;a9YC/d.,^27P6fK
&=N?X(JEUd.&Lb?MeaAC>I&e4OgcGe5:73Vg5d3ML>;b02=H>,?_0G1=ePWO:WL.
9[+?H,?N;LOV>91JBcO3[01X03.G#56EH#gGQCP^CR)R8?Y)NCS]ZE=Y9X,G]AHH
2LHUO0#.75[Y+&P>#)\(YV;9V>B73Qe]W;7^+HMY7_#-F3^a3b<TFBAHS^\8&7CU
gCSHCZ+IQN?:Q&A75f1][7)aT?&CgaBN:RO.<>Cd2:>e0KH)CP&P^W.V@YT,d>I8
>>.HZWfG?D(/_Ac-Z+aCa<[dD5e8094XMF5?J7^[7Sa@V2IF96WfRGO&;I3IHB0=
VJ)709K(5Q5gT,MCbUQ)IVKI^C@@:O)b\MV6P;U?_(3D<>HT9K+GfUJbg&#A+SEN
3(P?#E+<96K-#.aO2Wg_aWDQ>/6[&]+>HeH8G-Gd/AgJ)IR\eM2ZVQB-TRXeCP4=
:=][M2/RELL2F?GG7aD>619c8Td\^B)[#Q&f?/Q4bGK+bJ(5W>ZU&QEGFDa0@7XP
Y[SAHMIPS_g^N[U,MI-\[#3(UD1[#8N.3g:@V8U[[_E)_9TOLW[4U[e6&9W&F8H=
baL_#/#NRR<SQLfdCU?KKP303L;0]CUHJ_M8bZ7aeR@Q/<7RN.L<(>c&1HP7QC#\
1+_EDPOYeSc3#XKH&R?+acH@de-,XRFT/>HN]&+.S5B3\G2I85[PbP#<XRP/W@#N
9Q<,(\0,.Q).OBG_HC1>Z]1JW58F-[,A@B&X48/7PS#NC\B=\0H9b[1f(-D(H&(c
087SIAX_Xa];2gB]<6<EbIK8ga71DPFA(W^b?,)\N5?bABZ76LS+<9YZER.dAb<O
3[Re^?G&eAQ)/9/G.:U?^64fVA.+^#T.8+,[c-IOX65R]E:L=Jb6I[1&0FD\eP-S
&1[0@e1QM9XL=MR/JAHGI484,F;=FGURgTdIgG;.NaITN^-M0MXDfNdaA,2#:X]<
TP(EdGW7/)?;948NA/V2>Q4I+[a@H?+]2NPX_3D5#f_(39bdQNCQ<V@f_+=@/2+7
2e1=bd5O^9MC&FYLMJ?H0(UH^J:^/U.,E+&Rbe\bO<Z,Q>&GVXK#ZgdIUe>1SUa8
cW,9Q38(<dEN&a2g9=,N>ZT^b/F(YG5X=K.OO=HDBSJc#TON\5IIFV,S./(&SVD3
[RR#+WaMN/EEI+fX5+(D79:I@Fdg0EKS_YP.8OC.R;95YC2\XRNHL]DS6;CSG0e5
>[b>@-C4B]fRNWK=JJa&SE/bZK;3E.-P[c[_eS2ObR/<=,8/dQ&@481aRZ=EJ8bQ
Y=dME&=4RB.-F1L+V&->ZD\PdD/9NUOgV:)(4\,4UBe9TU)2bL5d,dU6)#HePS_G
BLC_c/WMGNOML[LL)#B9DbY]HQ[RPR:AMD)0QDC+I[CPeC10O4+8IRT2+:f[24\0
FPDT<ZB57dBH#9W3EG2@?P\\Q;65JfFJgJ[@NG5(9SDZY/MG<]57_1:Cb)I7OEM]
?=dXC9c)X6D<39;1Q63bO/-1IS3&O+Q9+[+D38WcfGH_BC_#XJCeAD&N.>UU0b<F
L/Je(6)3BT[e(<feEO?T7K+-60(V6;1(OA1dJBa.)3gL2^Gc,Lbf&fPPc143P-IW
<TX8O7F50T,H(+c>f\-;3_V,57g:bdI0C^1:KMH1\_5c06;V.6]F,a=9VN5.A.K\
Gf5AADM-cC4H-ce<7&]LWE<O1gc02I#:.>Z66X9VC&-WY/515d:SF&AgENF)fd^6
&DPJ[_&UY\Bg3;)IBeZ5Df1)b]KTac+8-6,&9Gb#9:,0-0?V2gK]d/K0fb:GN^/6
^GaW<Y=<8<+-9^?XL2eW,][1<(b^Z8,NOZTB4>0Mg_?H?),)5FQ6?45E&4&NX6?@
d,0:bGT6H4DZ=geYWQJ_+.Y;67JK#]A2Ic;)ZL0b5b,ZFQ@&b]V(\eUS^HOB;]9[
9X>P#VA0bXKXB@<T^X7[M8d>9(BTGa=(57C9\@?2-R^Q(LVY]YX8)</aD@A9+c\?
<5M6_R^=PFN9S=)+Q4)O2C=c8_RADRNIZP)BK-d^;QVP(Y[]2=U#+\K5g\)Fge1I
)1NIB[P0SWB[W=[b6<5_:IId53)A^b:aMKcPc>/#CIM7F=+UE&M,.Q-bA7aGA2XR
BH+&A3<VRgQdVE\9OE;@OI7GK4A,f7F)?U4+R,WB4?BdMc+30QHbH[+dCOT#WaY5
./+]H8Y_;KN6QW?ZQ0Se9XePKB,=Qb@I+82,8@K<bT24OK5?3UBPO\YO-L.&X][7
b@^\[XNHbES&NF<I4J4095DOQBG4^CLJ]WWAFUD2\H2C9-S;^X3V=+P:@.JgcI4E
&J9F,362;H(]@+R_G3O<8JOR@M3XcY4)bfEGY\XZ&XSH1J;[^b23_:UNAU6SX/Aa
DBDUY@WDB7Nf(/D_5XL;^6W.31_\EEa-[MQP2/HZ)[QSRR&eQ7WIGURc<M]GbU-H
5WJfdN-H+_QHb&a0[L1&/Z/A=&/#_cR-@8bM0(W@WLB1#aO8A&,X&:T?e7fGCVY-
.AN.)d0dacF&37>(g.\#Q#).XW/:N42,GKG,>&0;gTYPGEU@>f_2V&5:T=ZeG]31
N^WEKPB8L+dU-HY?=;e66#CZIP/a&dFe2WbH@M5;77@P2WK]SJHG(]gV)STUB(LX
d,F\W&#6cWdM(HP\a=9^V</US\TKK\]^GP;QbRNF2NJM^#EX6M<YMf[SPI_X-E?4
+DE<G3eD^,#JCZYIPLIH^F7EVZ<4FJ_-=PLFFO>9?Tg^fbEb.Lf/_Y2ZL:8OQ&:#
9AKY(2[OOP4(AELOH;I&K#FZTKAE3>.6IDfY1QD.f6GP5VZdMGU/C,A/5e]@IOOZ
8C-QUO7P93I9#g(1FM<7=CR2V12:EcL:N/=:/cT//0UH3^Aa<SU24gaJD?X9L[G1
_<71LgI4_,f?=eZG-LaDDPW^+Y-,DXY9,R/V4H=T8Z+)N;?DA+64NGDHE\/0KYMU
I6Tgf5@^9]?3E\2.&McC:QWGLR>DIe6W7[MAP0YEU\6-P/eHVga-CWPA/PL3YP.-
QMOEGZJ?)bQgD:M,9SH8e)3.b;R7&2e/FX:,[1D\Q2&HB&dQ&4PZ&]ON@+5g:B0E
?N,g^\KR<_CgFRgfDVSC4)MUM_A(0\Y+c[@D]E(M_#dGP9@gJ^a)5VD8QP0D>ZVK
MBO1=d+TV]:V<ScS9Z1><L::[O<H,(7)-B;PCa=^S]]2N)KJ[VX+b&F=6:O\O>4U
OSL/dD,.Nb_37?;7W[9S&.90.0-\YeTd#J7V^AY(#2>#1>8<8<0PJI=UcWQ91_VJ
YI1_eKGYC7G(X:gVf+6^ga^K@MY(-<dJT;/8N_b<XgX##CN?X&B[_FARG>OX2bNg
@@C[5#6?AQ,\V@:LQQ7Q<X&<1CH&J6KK63:J4R9@4K7&\^N3:DD>P,OP44TD3T-8
a[Bb(FJaSV(a;4U@FHQH>[FI<f]#7<]7&.>\cV8BYY-;QV]@#]\#0Uaf-\E\8&:V
0U6;AHBC35(9S&+5Fcg.R7TIeL;YRJ,CA2O#^6e/2EV82e;6S,JFbWFb63B^YD)Z
WXa1>OcAe-\A1N.RTf6)W>U#D5-5MScV(]@JH5ZMG.MXBL9dB\/JV?H]GR84<&T)
0)LQ_]DdFU,gW]0V;.YV+<XRFP,d]=LNg),ZGGEfC\NRP[.F?AB]eF]Qf_cJ&))X
AQMO4#<;E>).Z4<d7Q>ZJL@R49<(O4X@6G59acOH)b.MPFY@+b4#:^He>_W<?N05
\Q@?(+1)&T9,=_6BEE0VF^SXDG=-S+/:R8<QIcN0<7&:60->@O6_XZ=X9EI3+.2+
\QQV)Y@BN?f#0E-[4-DQ&XIPYWADFg7fLFH)>D3]0470OWdZCJQ<;B;)=F2P1JO8
CN^C7K?WAa<bCZa12G^/-3DZGLGP;,B<EW\IP49bD-c55<fOG<,Q(4OfeC-+@e3@
=Vc=OWP@N:XNa_ZRR/>H:?4VR^#M]_1T9OQGZ5QgQW@Y+3bEB;;:M1HZ@)D0[Le-
^2-9O\-ZU.:T?b@3[P9G)We]VX0A7KB8&,8;T_]U-Q6;;a#4La@AC^2U5^EUGA[<
4E3S34_\PFBU\B;J2b)_;=Y2#Ud2FgHVK-.\NdUEQ6\/FSPAGV\Z=UJMXf2U0]DF
);[<?UZ6W1X>P_6N4dRMPUQ,I(-6E<VS7IIE?>NR#bgBM,:TJO;DU+@:^Hg#/)&(
70AG[bfd<<G-T0<&B=&-\5)A2>=QLQR(&.AEN2MM,^\fINR4IYU,R37=TG,]B&5_
^222EO(L)V#6XBMR0A4[b4\Za.HDH2cf(T<b.-.\cAMacMJ@+U].;Z6O]7Y\G)0Q
#Q_60;YTg(@T0DN<1YYGYdV/QX)V@bZE<K,2.;K0&U;&<SN1<0LSdT/D(=;KP7;&
M(/Mfg1=3[6;cEF+f[EL^]d:Mc.JHfbS,MJQK-IZGS\8.S<_[N/O6g/^>YUQfU5,
X:E]_0\T<A-=)OR.W#]1C&SZ+LG#.0;FNaB]cYIE<Y4)aMd\#,,05\ZG,J?S<A]-
]^5#g)gV42]^\97<+#H^d2L81aVBe<Y2F.JQ1FP#>LN/OC<ZO1e12(1Q0bB8e2J,
<]Y-ZZe0E/e6O&)MDY[0\a8[0-3#?9IJBM+3RW/164<XN(6d:B7]++MCX,&D5@JA
>)S8XF0=3XAGF/d_I[^5S)I\KQf:=a>8H8Y_T=K=N7#^-RX2&X;6WfT\#D2B5+@J
U6++,1X1[&-fMe5Q6aMEAB<:@Ag&]V,_P52N=-cEefgVRHcOJG&(JGWZC]cDCaT#
[^_#G<LdH[e;)Z]#YU7<(.M>SUG>4NE\0-04fcO)9QQ(8?)#HL@IBE.MRY6:HL];
@:(O6NWcMU)IBg\^MXXfXA/NY^GCc8_Q?RG2b(KRS[:TUWF&+:3[2]&9-d&7Q]2Y
N/L0A]>MLC\GZ4[M7@(C]g3)[LM5#^8c>Z,K1a^EAgPC+5/FR=5V55TW^Je-[d:;
NfT2S#;<NbeF)K?7_;-&f.=V.TNW#9&3AF(OVG53g?^R,\]J7&:NHC63^.79__01
Q&6a1#6MDdYOK815.5f,c0)\9L]a(/;g4PFXC>)+-+NMe@:1VF(J3aX5(/Z)Z^OU
+,POSDK@UaaQe_:a5PcUQc:OX8PG+?+UQI7Y\AdbKTZQLYeb@c&c?A1F^SC5B._,
6F,:M]CG[QU<]LB=6+Ha.PML,7KV,g@6a&,)6&=.@g+2DQ-\(5:N=[&SV?V6L+R1
?.ZSXKCEeLS.ISWAF,AD@Lc=++a2Y3T4?Og#eWH90Ef\Eg6ae=E63Bg&f6Na7NZV
&5/Ke0DBB>BgO46,JUYC;cW@9bM7..49e:U(g?J-1@c:U#[O9)HTTdC@/9/D\)H@
:,PX2TQ87BCTQ;]g+P9C,)23E>D7>/+<A&@GDJaT_F/M[_@9WEYM[NM/08BeGg<-
=2FUGPO]M?I(FfH.1ESA)M^HT(Y7a6?K;4U<CEWJ-],48eDC1g]1DBK#GbCW@.[V
I:\-7V7&#+Wc-S_:AN4=^d48^+SL>[:J#,N#\^BAP>\bJ7=DE[DT]GQQgVI\L[C/
+#b77N<QWZ&(T.#fD9ICA+b[Cc0b^D\dM3JCa2(6&+\GK+ef9_F/SU&+d,O?e./:
gLJ=JZb1BSGUXUZ;b&TR/CW?.bb4)5?_AXM-N\H\,(5gQ2N>82BZ&I8Kb.7)\Hb(
b7KH6]Z-G35:14<[]G_Z#.1U\WC3;AZ2/@?5F#e(R@.<7Q&UgMC27<0gLE;W-K/H
G(B9+I_[=&?_.(SNSe_WV,PV<7d4F2-?EF-C^(b/1Sg8LI3@D_#LX0e4FC-3fU,_
6HGSV;5O5IH3O61X?d6O=YEgaV@Q&_BU,e6[.b2e(C/f6+CA)/48+MA8/Y>>ORLc
,eY-+KD>TLQT9W17B40NXM_2K_Q-GC3OdMOIbVD#-(,WD4a(@>N;;05AZc.V/?;)
HCI.G4\:H&GFEP=LIKR-\L&IP_K@M)RgB=#?O;2=JUFA5G+LO^#bce>]@-V2W&Pe
GS33>)Z<.I#S=:_,aZDZ41,92+7Z6EZBBV_1L:QVIP\=c6\=\dHL5SFCEG,2dFCI
\^&b0;3-L?DF>Z7,X,5SPMG7ed.#)+ddG,17.b[>OAbC1^B[Qaa)EFQ1HA/@RVaO
M5&6EaQ+0V?<IU>U-dN1U)_U6g<5)V<XVD5ZDLJaJfLfYaD2YT#<0dIRb7)K><R]
I]:QKA,L>L3Fb[#F,6I0C<[BM313_dV-^_<+[O@=):c+g-)D@Aa]bbLeAN.(?&f+
QIaR_?JPR<@?JebBY>Fg-3+Z.1OCWc@Xb,f@^_bT;OA)J0=,52]e\2=.)LWRad@I
&?8^2D-Gc@,]c98?UUXWK\@_@-eGVT\0^?:U&Ia[==fF2d&:Md>,9]<Mabf\gMPU
Y]a)^c0CMGE55T@V1d8[(W\fZ7;cK[1)B0S_W]cdW\]FXIJ??VU870I/.)9J&IL6
@DM;b_IOK-IKP[:KX_7TT./Xc9U5e5dbJHN26MfcOJg^FAe\]gR#cf<[2aD\BR35
#Q_7TLFTU4b)[caQ5C=Y]X:NaI-FV;ae]NS=BL+e[0UOfD/UTTLcg/D/UO.5eZO,
aJE>[[B/#F<4PfTV6EY<._=.P0d.4XF\>W](<e_-[O]T-LX)+9W3JL2/<;/Zf7[<
BV==F/WU1\N;:b&Z]:1?g-\\@d2)LZMVTXHcR#:dL:]S@1,2&BQ6b=a?=Ne1M]B<
@Fd.^:JBR6I6fWRSXb^[Kg4a,JPNB)=Y[X(;CP1OZSH5Z2R)0gd4R?3aEE-gC6PF
U/S4[]]WA]5=PB<QJd2bBH22FM/DX3VAd-^MJUfQJ+<#\O&#;[(8M6MPfO8HZ\e]
G1;0fM;6]ZHJN6#/9SS/K?J<3H?SV6CF=-g-)0eJc1I,C&>Mf?S_gB.<Z:Z5X;c_
\SC358JNK1G3+J<Fc6SPDeP/3TJ<W;+]7T_L]^]5DO);KJFS7b+O5eJ&#6dg<<6H
/+cgWEQa3O=+=49a>A<@Ge]GAYU4]66<R0:SI:K^^2RAb1]9VP(+W8_XH<W]NL,P
6R_W4F\3#>BF-ZVCUEKIf8<aYg:bc&2G)\78a4N=74AaYXT/MF^^.fW+_A&;Yd]=
(R+Gb;@-0UR<eEg?:D\Eb)a<],;7>_8H+gI<R46S,6:.B)UfJ.1e=K?.K^P;:@V.
Yf^Yed4;)S?=\)bAQa3AN8T=)BNX4UAU6_b11JbQ)adMgV03/N?2S?T/01RXbfaN
T@_bC8^2e\2K;TgAG(3T]<GJD2d#f].AL8GZ_N76]GDg?^g]^Y:@6fcWAOTN^@:]
O4LG;8:66bALae]<P7TO&W@VgDAV8\FIb;aY;.^@JegY[^fCfg,_;0MX?HH4(GZ<
[cIfE84Z#-Pd[g8TS\H3U=-9;42g]AFe?8711>a;J_GAcRW8)>NC+2?F05RFP@#_
]J4IeGLI5S.>9WF>0#&.0)GO[:M\8A,#9OZ(O=.MBa[=dL+g)0A,^f(g6E<9>2Z_
?QSR#Z&95(@;)[K<+8^<0P?&>IecY2+K>X+<ea=H]?E&40MPJ#gPeQ4Y-#WA+f<K
<,H1)g>KU<b286BHaO))J@K5Z7RI_e,FWE^UQ0B(.+M^F^)BDP4J64G7;Y+L@PB?
Z^O8f4F5:d?1FN[P-7ZK[IVaU\M1RbQIKb;/PT.@V[2.S)<Y7>_Z(-+J]+WQX62:
VYgYB\O0eTT_-[c]U3:7/C=QP?6R)TO3FRACV@]I_J=:K@>F1+4,[:cG#1=EL_3P
2&=Ha7_bdVO31]X3Cd>FWSbE=b/&[PGBI>>C2Y9W>;BZ?7[.4+)adG1I9?+N8RZ=
I-CC3;3c3>Rb\=Fd[cE?1J_6c(>X)bPf1//#&fP1)K9VQYG3O1CIa[_@N21g?-AR
[#7Df6O:/+@Q85TNQQ?+YD(?<5@8_<71L.T8O;_Yg^Ua9+=6cBAc:YI#60:)_L6G
0#E]3#T-F:a/FDcMb,Y92:95-A<KVS@&:]-Y[^B=P&\_R+FJ@@>LNTV;[V3[QK)a
S?DZBN&GcdKEAU8POd84I,C818C:0HcgD^P@\6Oc[ROc8a:Ag\;J&T+b[)-fbW9#
L=(:)AI,:8PVdE^>DbRCJ_J9P[e6Eg5L_^<bBLW@E:GLR7Be,FEAg5E0IF98?CRC
<E;?:S4H9/U,K+)G7R.U=]@BRG#)gBgX8>^a79^dI8-ed,VY0IYW+GDdEN38)T(K
0XT#5K7D;<GGKe??\0O,&E6#9g[1TTZ0<,Hd=R/XgTHIW,-eCJR(0F(?A(C7-LH;
Z/C_)Y]4NZEKP4A4&WENXH6H7MAH70^Ic/32XU+_+G;T(S^+&G0#3CHc=3G(03Q]
=b:)=4US8Ice[R(gH524VV#)1gg50=N8HaWbMIA<:gQJ5dX_VH,54\TWb)+BIS)]
\FJcP\\TEP-CEZPHI9<:SRK3\S36FHP,Y>\T<d4?c;2JAY13TF9]?U43&-\d=5[5
?I_1^75TVfS;(8RFFS(YHVY-K;F);d47NU+CK].\A;+^V)P\C>E?Q;_V<)6?N/gD
V>\,:80fH[bGceY,S[YNJ(g289\b3ffD=A=.8):)CXd[1QGaUO.(87>6[;ZRA3c9
bD1N<-Oe/EAQ--/TC-?HfN9H8]@N9=>Uc9]@6CKKL</>egec[gK_<_a+N@12)V&M
QSg79b3dbUde=PXHfNgT(J1EK#UJFLHJCX/)I3?fQ+aeDc)dLFJUUMN50#7]9<)U
6\ZN81IKR8BJFJVBdG7?-9ga[?&1ae.eD7RVQ4<2J6;47;D[3cWgD7DcKJH1#WaJ
P1I6#:+aV6cc(TI#NC:TNST(FCA=22NG5TE4PIb@)4EW]7V\aeD9V/JdAcB4Ra>5
IX;W7:UH_G&DR6/B>)P:W]Z2Cb+A[_2^)W;&UP)=2QBdQKaRCR.db(?POTF]b)/f
(0?,b&&S@B3K+3dC<_8C105>NK916&?M&0TR4cT-[cC\98Zdg-+6cI;CD>E034+#
X^W^Rc#F93Y=ZDZR_4_-+K5O0[;N+2[]?>11\JH(89T./782/+P(_W4eHST>&1D+
^@KI_03IKJS:+R5VcagTF\FC</1GU.3OKI^9YDY+?4#+Q0#5Hd#M;^,BRIU>JL[&
5]I:V^4D1FYZ=aIN1>):F:C4Y]4eG[7;F8G]Fe6C\\H23cY^BO_\W7g[L:.+YQ38
cMgS+CP\2)U.17/UQQIV@WcP^?FF6<+>B2]5B[NbE[+Q395cR_>AcC_8KS95CdWW
]P,CFC1T@0dKeK?NdG8MPcRML_[E.MT]S<;Y4V8bZVQ?g>COgEgHe-U9QL@4<.Da
>_fX+DPKOU2(NfU=WH<;GX_L3a5Z_/[87L4NREE+[#OgML@\eLRE8,[<)[=HS\/<
<LW#8E#H:d+<XGDC8S17a9Zb:WfTTI4H=4OKC3P(B[1/g;?d[WcJG;BcK6^TDgTF
8L7[,_5MVY/Sc<)[5Md2);YMfPT_57&CPdP;c@D<]CNA3Z1YR6G4a.3CTcF\3^JI
8.(5]5S)(A+T(4ES1YQ=b/dNYVX/XZ]C8;4NA5@D2_dOX[WYK>41U7QYA/e[TgS9
D-RO0_4,dKJNf?_>(beX))[a81.CFTQ7/;^5@2O(fbR65eB-(9C?,B:XVJBM/gLb
H>4f_V?-:S2S2EbMa5\=Sg9ON8Z931.HHUMY7c\FZF4LLZZ/(GC&B>[-QOP[TH=.
68_(X<X1@/U=RH?T:Ae2f+HK1=:SJN9bOf<:7KRED:e+^EH8GaC1/H<ZMQMU@LV/
QV#=K8-ND+Ag2XW>,.9e)>+@=&\dD_>dIVG^6DVEE^U[TWC8R77Q?+gO:)B&Wb&A
eXSH\8eAG8.9gB9eCI:E.5fJD>UUCN=aGe[-L8/Q@/OS2V&75CD.YR2>#;/@2)M+
WLVDf\ST_&+28ZX;T(aEANU1V;5[e/5>QEXbQQ^\I19SV&^gO-=QGC6=P7^I3HF6
;@\cZY2<J)N)O62NI]C6a^N-c?\=N9I/0M)]RSD[eLZR0&BGg2TS0d,7N)1/4&a[
T9D;@WE())\?,O99V#^)8JeY)J.3(0D5;\<aR.NJGU4QK(+VRNRQWOG&I0<a_C=S
7Q)/#,285OO.>Z#(Y@(B/C&:1]JGPF=.:.&=N;)aef(BIQ)H:6gfb4Q9V)UZ9_9g
]JX3eW\T?Z2#U?[3X^7a>,QePGf^;,Vaf2_T]d4>X;g;gf9Mg(VR?8XE[<&12Sc4
S1=]<P[CZB0[PH;4B/?dBYO_S91&J[Bg=?96#L0;I/Xg^)VD)4;6g63A)QJ/)<I1
D;@A-WdRJ8HJ483DNA/L:d]a_<b=#T,N6U#2dfEA,^IaG[#.CQ_));A3Ve^:Y9f]
aV(^<<7RJ2O4d(#RWZD,KY>E8HWTFIXbWaG;XRV:[EWG18P#F@>6&DR/^<_>AI(-
(-/,60[L@E4LC5c>.VSa&e#5FEML6@^&SaBK<[YFAB44L9PJP7<QN?[]E&M]e<d2
+,^9G#C(Ye/]>GIdD5+dBP9L+;?aI.JFC/D[Gd.8(,@ee0,M^1LOSPD)HFf&A:K4
d+K4/\7R7X41]ACf5J1c8SPgRXbJ2I&12e+[_7Lb^c\=P,PgL73O_6T5gA-+5L3C
)T<,ef<b<8>OEIb^/g&Fb&Sa#HOT52#>32/3W]b3Uefe5]8_&KWf56Z-1^BZE5&M
/T<?a+TAI+ZcCD.WP#\(cfB)AH2\>EN)N=_-ZGGVgeICeFUd]:,JY^D]<[AVE_<N
a2U6fT\gACdd\c>JC&:MP#Tb@B1[7Y[0[D.2bV2.F>],N6M.f)Ib<dAZUQ[([b/.
.@H3G-eZ3;TK4SIE4GO-+TI3?^.(V]e=Q9883L.E(B0X894@^=dJId(ggBT\UYeg
QS?]cE\V<06/9K1GNg1I4GRRD/gIC\KY@3QCDdF^K)R8G0FMLJFG#XF?UNf[17GB
.<e6^;3AaL3S+<O)JLH8>?LDe8G8]_029<dRg,b.0Vf#()7A(gcA::YT<0Zbf>KJ
[597eb].AMdd6GA>J^/(<,<8\;Z<E.YL<5B+d2X/b3d9T3N2I/Qe3Pg,X=@+J8WO
:eB@a)F]2O5;:VG=9e+<:KC6<dB:M14OR5]#N\>gAF/7<KPN>2_XN;V;G^a5]^^\
+.5TM9XT]RbL.9:M5BAGP0(+JY(86NX=OHgaD3/2C/IY@\P_>EHeUY+gF]8?SFN3
c1E>ZcW=8OQ)PJgBf\1>6cB8e7Z6FD2R:CCEg])cE6\.C_,]^Td0D^-H/W:BRa+N
&;,Oc>XT2-KBTAB1;-EJ;C?,SC[8Keb82a1eaeXP@?]RO]L(]G\bFIa8]]57D4GA
Q=7X+bb=E>F\c3MFd4E->B4XT4L;S=BHNVD>)c4f99HdG\0f8/Rd0P\R4cb9G_?Q
.G+=ZG9?R2^+Z:,(#1L].+?>CNV9cY_^B+ES^b5Y0._G5f/NIUEc3HJQQ<Q/a;IB
>;M1(aARFZ4fCMJfVPg;1S4LYRc-.X-OK;&GaS\Q1aB#fV8dM+N0RS_L(SN;D-ER
fdbSHbCgAR(R+[ePg,GP0gYUM([NX\I0IR>caD/,DPS@=#6H^b/[Q/7+<<8\-Y<N
KJe6Zd6eV,9LKgY)1gBD80Y=:YRX.;,OcZcR&&)L_Y8a?/Z17R5dCP]e&=a]&MS<
SXV-MORR=AVBB\RcYMY0DTE@3Sc<2_5]I_geYd6&_(<?G@;\[LC+2X0faX-R+M-C
E31I9MZB(T<T]U+VU;8B8BcP#X#.:,PPPP,gR#/6=UJ9E@.#[a+/a4;4GbDOY(V4
K0Id&B+79TJHK,g>PeU4I5_=5\CfG8VY89OdDP.Z&?KCZFIH4>_VR#H)I)4c\VWf
03ad0G1-#A0EBRUD286[IB,5E4@BUegAONN#,UeA.LSIb^:^B11fd7IGd7&BMQ_^
gLQP0Y.-5DPAd2+b+J5L>dbE&?Y.]LaNA&/^E<ZfB,Lae5(X6EJR>AdR]FFH\->R
S)T3dGd^E:?<D:?NQDY?SRc1aD-^M6^3c_L&CG;T9-3g4YTY3P2@bQT_<N#/B02B
=<WggRO:eJaaB22aae:Kc+.5.7VKAcLVM]P17CO8-ObD/=X@218X@G#@POa>HAPA
T[HCWGC2Ae;1g=3V0ERb#16g<?&,afe6d&CT7-0:E[:R3N/@[O-_5PTe&U>@N@/B
D0=&RS(.9P-(/\&+H5WcZ+=70N^bF>-Xb;F&1GVaG)@I)eH5+MWOAI)6]Q9ce;RC
BNF8^fVH>(C/#MIN.Y+2<Mc#Og-=]dfP^)(M.HM(>TOXS,W(NeOS2<7P^;Y^?];_
SIRU;28472Q>L8,W#TBIgU_:HeT0_I7H@:^;:7;S5?310Id=Y<DUR[.aa4QN;&@5
;&DQc3a[X^Yf?S0Ra8V3WF5HRG2-8>,V463&?[cZPC=Y+>=4_Ye,T82F0S@Z&7gQ
8[ZG:R/<K-1?=^I&<U<A8<33<;g+\A:F/6Q\B4>>[J2DLe<3C5H)4[JCP0(ce0+?
,6E092=>YHWS&N,,^IXP9)bOf5CV.]E)?V\(92G=?>\<bTA.Wea;GR0>OL4VQ@O=
P&U=e1\+324dI>@UGAe8VSRTdP99?-9Fa^>HI,U79@V,LI.4UN]A8/RBTd&e1Hd^
f^<?,D4MEC+?1Gf]IacT)A@VM@?R,0BMF/LR]fX#<FKc5gGV<801QC@.fWeUb(/3
S\@/MOE#\GCPZ-47[+;ObVaJDV9^@VRLGI_H8NO],E&@.S.;d5W3)8-O9fQGVSVf
He)UV@8U9GCWg;BC4c&gHE4Y#1-L4IBH5V-=C>]Q;E62Qa5_)GQ@\F]L4A4SZK^g
C8:EbQ/Z&;)NW=_55O?-<fRWf4>Z(P#@154M2LF8Y/\Jf6PW+;#S]B50cU,E@:[(
0Be+B)g<,_GB-M\:P5IcNRa#Y=\Jdc<BOV+Oa]b2.TZ7EZ2&O\IZ9MC4K(fAdg(b
RM+;C\9a_@I@4QADF[(NW\:-;+;3;;OZHYQ(&aW7QN#CdSH,\a<F<#1Jf6>U.g:[
7;GHKL1YNY,F(d[geaCOH:M.e7aB(FO):GJXeW>96[/Mb/?NY60(6?TN994/?RSG
YN.f)M-TI2X&AA?L;?g0(VTd_)(.f:4b7JXG>gXF9\3fE-TY;2,+EIA/FM^Y>3XZ
3E32QR3B_ZSJE1,C3.O_KOWF<IRJ_.=HJ4JPD)TZ:66a.M&M/)#FgBUTBL4:W7?S
S.=D&)[WN\Aa07B(D^8(7V5T;\41VcBES=HD+35<[f\(HWJeQH.O;-HO3;=+:&P]
d3L+<KI9ARbE0)g?C/SD](3I2DK[]HK5KQf\5gH>C9b[=[Lc:_X;G^,6UfJEIWWV
T;3^NT(.aOB/8<DZL^)V8eRC<OC.T=0)1+U_I>P>7=Y:N4W-eCVYUJ.X\DYR97b/
a;=D+OC@Y4N),8+L<_0Y#<dQG@-HYg;.F@16P+JOB.:G/FSAD)YZB6B<aeMH23\A
f>T9)/6?d_e2N6,]53Z/_@7<&.GM])bEg^aYdZS8BJLdSAKLAJ.#<CAARLBF-+d7
2?=U@H<I)PH.88@=1L,>R)A]1T-33\0NV(#FRM6GT3U<X.<Y=IdB>#U:;U7O1-)Z
9[Ha^UDJ7NVSRXX\20WfM=OEXRd]Hd2AH?M[.Db0//b4Ve3d?V5EY0TC<P]8E7)N
IKIUaI,[SdPGRSLcUK.R^-N;d=@S+/V<A<J:FPEO&;+ZNX,=C92-:#.KR?F128MY
TQ=QGTBa:INZ&[H47K2XML[A<R(XOb5M&?SD+VZ581+Q)2M=\5H8CX#1&+?-+;A(
Y\d&.5L-5UW_Ed>Z_\H11VBTO4Ge5Jg.WWCb,ZNFe:4:gTJG[TH44SXRCVT\.@@Z
,^OV/_39T#c+\Y=ITM309JBJ;^&Ve8(\@)J=\;9Q0bWW2R0DO\G91X,I&M6bO094
HP:_9=@Ifg+LKA1Q54DB_2]a7>\VP83J:a)MOKO<32?/IRVc<;=aW>X>f_S9M8ad
)aG2/RAU^a?.J:CS-a.OV.I>>[>76&bBEg2<La:==>A)d\_5BNJd8KXec:Ad9GIe
QJCI@U,JX_#d7>JbJa@+&G(3HKb\BI>)]f;KeC]S-.B#JMIZ[0ePZS?fX#&[7WBQ
,Z7#8[/g;8D0fYf#-cQ4H#3^FBZH#bR\Z9eC@dEJ6C:+P1?2(LbXd-Z9bA&&D;^=
@P(8G88/DJ@O?G-B<;W;Q(DJbB3WWXfWIKDYU3,f=3[1DD#6.23GbO#SeFDU6[>L
eJU1K?\)W;6b>(BRY5P?G=S+=1[27?WE,R<8.cU/KLQ2\6He.9)7<TKBLAbHR&^)
]@PR,b(c[@PXf2bDF3TfCQ\c<2HL=CK(A&,UY&dH;BL&fC#4Pg/2VMR7C/9@E@E[
[L6c]^Z5DC(0^PY_AK((_1S1IU.#E;U)IJ&8_7<,(,1<(ZX7<T9@FV.-X2460HV8
@HY@Af]_P843ddFg>ZMQWLeOW(C-@F0A92G,UcR(d3JaP;VTTK5+O1?;DJ\H>J/d
N1e&CFe2[<9L3Kc#0f2(L.I?&TDPQ>.Y4K^#TB84HMS.^UMC&MeAAc3#5F&\FRBQ
K(TBAa].5:@UeJ\/Y:,\RDGR1ZII>dJG[d-_b.H(5<1KO2Q1B/O/.FELQQ/O/:8L
7dHQc[.4NO8&1_13aAf3Jc+F)X]fg[>CPSVIL\bK/<;8U+SED&O<f_PeXQ=>E;G4
0#SKLg&424/U=S.FeJCIZLUVTX0TVdbUPd&UBf@.53(T+.a,SeW^PfQVLIb#1.T-
Q:bAfNca\_#6(YCTSAR+4IUaNBOJ>UMWGdc78MI1>S^+2Zd#)+)dAEB,>MJZC4H9
,CFfZ6J0+RcJ2?Lc9-LAR(#]2Mg0CSY,>eN@)>/Sd1UBNP[ZMM0=<ZN\=9H@=U7?
1XEDg_=1P5Bf]]4735e#SaJUf\JM<S;QM1^@fcW.Q@gb2eLN,;XGLa&<A(5gPGe+
fGJL@[BYK9eL@OT085WO)U8TSd3DdgQY14fZecPAR(JXFEACQF]QVAOR55B<56<U
E62BS@UI114A1PEX-8-Z</RBU#RU_TA?U6aU9^Z1N<b@PK[[NO1O\b@I,MB.RMd3
TA[HAO0DZ/@:ba2Z;,N<ZgW4.1/MKG9.fCSJT3DKRG:EbC]R];8+)fJWe9[8E=SL
?X[6;XY;R4_DF6RP\37DUeGB@^ZUXQ4AD]H/e_)./W2/JD4V;V[OIe6E?]5X@3G^
W-PX9AEd1Y6_LK1J&@-U-53b\L\F[MgaW;1ZbX1cL.72#0&8e4LM][IDCe?)bRV)
RU4=/8#(>2bV<^5gNK8AW0[S/N;aM[]VbXWU^+WE#f=080AJ8aJ\K16>P)B80Q@(
LR.6?W5aM>aBTH/Xa99Z12S)@B]N\-e,H-,7W)G&U[O>W71[D[<&<b0]c2NLKEd1
B-E(ME&-@WIa.-E:Ug0L@OF>J#;,8N(,Z+<-6:RNSW/T-?R8Hg@^(5X_OC0FcgJ^
fR48T<RgE_)\7PY^JM<g\-;_;F;;X9F52PNL,#N:eQIeJ1;U#AR<5bG4=GV.VBa6
b?Nb27NeMW(XIZ>9PVF2KX8=X7TY8@N54E]AV<3L@8F^)&]OLgS@MIbf8&8N4AJ@
18\a@;MUBF>8cA=S.?R^YMBGRDEC(fP5QJK4cZ@;ePLcUA>c\KIU21QI&e)6abNE
8[LT:agSN<1VW>^_D1E=B;d7#[cYH2AYL(+aA,YJ/OSV\IOF/gQe#(NB3>#:D[[B
D>?92Wf(4&O<VReP@83\SQ5aKC\Y#0-),P]c:)N)X)3L+18V&7Je5H8@A\11E@7+
e4BASXa2:3+d&L^QP.WFCLeW7>W,b&YQFG#^,L>+03g9BL_XNKe^)-DRbeN^OA#E
U;)X39>4E,(0#3(gE_]c?0RTDdW^UYV<W8>f;4C0R::9MI57.LR:P[)fZ\_=AS/K
dLT/A])Z:IF#OcLZ=UC6\(H:1R&@_bP,MR\\RJR.A#?5,gF>fBEVA?-QPKg3dRa6
_BQe9MWDU@3\G)NXaF-IO?>3DT7BO2:2XPHaN4LPEG:DN3X4I.<HMgDG&,_BABT(
=>#Y]V-7DSLFM+;#:G70H72C.3?L;/URRJ\.cQ4OH^RaKN4caTNL0:^]WLVZK1:(
^JW/+/#P/;I@U>X@RII1O<]^KQ+3NeE7V5X]/,NH)gdg&3EYV@d8C[@1X/>]YDBY
bg;4E(H+_[,N^;GOXE)@CV>+C^X_<I4/+;f^(gKG)ENUgPZ]@-(D14a2\=>eg?4W
@0(EdC;#.FT#0b^AU9_Lf2K8G3-JaYE34Q+a>e0NIb:QZQ&gfaf?<e9HJG33IPW-
K410LEL80\HW\V;2YK@6&+)7Wg&,d8Q<H7P/7<8K3G_L@J&P#N@V#dI:Kf16?M5Q
2LUH\\3<-SQV+VFH&PDX5X@?5\eI:TD_MIDD4e+8RQFY\(\M,QRD85N&aSeOQ:eR
>a4CS4QRd_79MQ-bCQ=F@d,SU4AQ^K^<7Qc:X,<Q^XZ00a@TC.:fZO/F4;&DO]7=
YSLC[4/OY>G[GEJB:dc-Q8.U-(E1\E[HKU_3AeW91(>eKSfIPdL4H[+:D4Z2KK]I
T)//60Y,NHY\AAW>gWa.SOdLeT6N_/+N?[GS^LQ(HTHgcXJBUcf4eeKVJ3GMVb/[
=;->d@VZZH4H4^3MX#)\aOcI[<(E&88?4R:&6caCR.aPCDb>^I:@TWdW0U)Rdf@/
RVP>fK#(BO.EPFMZdbf)^<ad6XQ=H2.YYQZ]GLUdgPNI)U,gNX8@b@ELVK-(ZJ4^
G/J^CZIe+F.(f7FP:+<->UH-a,7O_G2;1/.J[OT&AEZR))f>(S+TJW;J?3A<#,.+
4C9\MJ75A6PD9SKdV/7fX3GKJ.L45KcN4+O#3C]0LK7G7GSHF@7O85d)>9\L/4Z_
dKdTaK:LZQ)MM>f792]#YQ,UC^.6S-I6fZ#0U1SH_I^3f]dALYK_B3Yb9F>&^//-
@7VP-:@:PL3A:A/9DY4b23_9)(c3(8X2RMSLKJZE:#KdfVM97MO::,][N:36JeM^
;?T4eQVcJf;/8CC&(7HY>^;^3N1N\RRVV??80:6^&9)M__=>AAKBRCN0\629_F\9
IO3/XCPa2F^>?&^08fcRYYMKcKa[MXdI^=B:,HAeMOd+84<=<U,e:f1]:KBZ]IWK
)#YUHS2MW(&PW]b;P29,EHARe<8>\>aU/-/;9P6B)g:T9&/a:MGPWO]Z6UDQa[Mg
E(FX1b?RW@U>XLBIf]/,eJ\0V8H(U];)CWCeOV2[4GcS(d2:2[Igc0#-28ED.KLC
cR^WW#V/,K4WKGD8XYMe,PUJF\S)O(:M[S;PccPX,d&dBB53F^/UEY/=,RV,0Q-_
ASC;T12W.96]XL=CYDM2W^\.e:;7O+S[-A4+LP97F[\1H\8HZFI[<#\JMHLZ7/=M
\UKYg44[)1S:cWZ,[Q,JB7ST]V=;#ZE;LX6J_@NcV\.7c<XVNS]2ZW:&1W#+^C(5
IR_NeW2)EN/(<--fK#T74b^H;+]+>].UEa=>8EQ;373bC]6CJc)9B.0d3G7G&\)2
5YF4MT31M;SV^&<W-=0.9gR4Y5/U991-T5g?SVT_g0HIZaOK2_d/WADe(X)aF^1.
(]UV7?O@<ELP1aNSIdB9-_]CO5a9X;2Le0dAaf8TL7D]Y)A&,g&MG>[K8/MACVV[
bG7IEfD)SM+e@,1GG]AXPSK1XV6cIED(<?cDfMR9bJ_>f+W6+5Z@@?0eK#@4W^+B
<H,5@V\cgU(/W2fP:3FDd(USM@@-F+\JUY=9L,M0EJ4f]HZM269fQFQT>/B0:T-b
,2[_Qb7Q6WH25\^W=JJR+&5IX?);\J-E6^>PG-@JR^@)_Rb^3[_GCN^\=1X&fSfA
X:WL#EL4-1\8MTd>3&Y<b]K@FSL^NHL:>6J,-?5F?)N2C-_aX_&(V8Q=HK=QO/G1
8C#QLH.[(f?YFHLa4&aN.,W?-\6D#7#d^=4WcS1FH9R]>,b#8?DS16U5V5f7/FW=
4=7Z@M^.b;V#P/0)a9bJ(LOT=>dG<Sd5#HQGc:M8QL.d>0F6.;-ZT:03fL+.Ab7R
5DY7:W>[RV&[aS[I5\bG\E?ES<X.5;dY9UZ:9J+74(f>+-KbgfcI&6.P:M;f=dYa
b7/(NKQ\06(g/6eeQN4YM67P+3VS(1:B]NGF\JH@.)0WSU1CCZFNfgWSI]6=)+R]
H\^G;E^#Y,ABdK0=Xb^D\gT/68=GRMaI:HYHE1/N@)+3-b:;:1R9gDWK:/d?]Z6Y
/U4+.[4RDNS<)\5^PC-SXaE,[1O>dHT^/>f6d_A5>513N12.X^afU2#^Z.X7E>YO
@M/HP:CVVE+L>XW=,]U,>/W/_+e-a?f]Hg\59SK+D786/#deH)E=T(73e4.2g4-]
N0dU67gL2cD4bNK=?bTRGA]XbG#YYQ)8YA=Jg@NZ.1T4SS.S1+?C&YAO65&ALY:^
.IU^^;MF+?ZVg&XP:/9UKCQ&P/90Y^N>B(=9R<3I<B[?78.FW+7GdadM.Y,6/5<3
\2R;?7[R(E56N-,SJI]5F&.cH=N2K>,d[812RDGId,/@<=(LPVWeNT6[VL5SDd1S
&DQ(dXNfI^1P@CBC5RcH?#6;fgA6U3MO2R<?F_g3a-6C[RQRPMGBf1eb[3_b4e]@
HS31G)TVPe-cFUKU74XF<E7;Ea.X3U0IFQ/R.-AU)21e4I]C=)(7:H-6@Xd0L1R,
&UMf5cHJ5,fa8C3^)O_E5Td^K-AEWXJe0D8gYR(4V\+dgCS]]DT9UO1(bMDLaXO1
QCf+G+gS(5M7/)-,M2ALaEO,E,bH5,D5+A/WM?GHf+L,+EeP9^.]&TE\;KMN@=/5
Z4YOF29YV>MOc>e&FI(ZXSBG?SL#W5[RbFg9@aOgEY<<gN(D_J.&O1.BFR-AU)[W
9HJT]c@A[fUMVWT=V-b9E3a\FSQSY0U\\7<VG@eV^,.2QGYZdaU(#YA7)F^OA:?C
4?&(^V:CaR?;>5)e2eHVG\380IeA]^E6M7X;a[RIDFUKZ;a[/d^MB7)B-ANfNf6Q
b,CMeQYUS[&X#K7.DPbIUaF-DfHXc?=@6I3+/+a4/K=ZY8B0OQXF>[:JDfC2]Nb8
/0YeMQ\UYSQLe^/G7\+ZU0>/<23L(7-LP.]+VO<7LHP/gVgM^1@+R0#bLgKN[a93
bcT>A>)/QPgYVS[Z[XX0[2X7b5fQb2,#4+(,;S)&^Feg&I,;@;^LF\.C?.Z.;U_b
+)fX.)b:^>5(:D#>]HD-G?.72QZOaC=_PK8R(/;0QX:;Y6c=A1ND/0c=U@^1eI(.
bKdadH_3>].&c>&:C.^N0EFR;#dfJ8RO<PGdgf99_0JDbPDY[4LU<X;]G2Ib5Z@Y
FF?)61AV_g).,JF1T,TO>>3OdJ8B+80P(@5T&_:)S59<::]K0@15HUDX:QF<QH]9
D6:6O3.3]EDZ.8A><XY#C_:)9&^B7OS<TEHE^#S,9Q&.#JXV3.)E(DYW^Rf,aKQe
\#1_[,G<8\fB.CSEc?38DCSDgfFN4JcbA_YSW\-#P#Z0UE6dOA-f;&d6+U>JAfaZ
5/6;NV&_,C->a5J6dXE/_VL=0NVb?X1gJF_B&Y1e4Fc4).Fd]?+2,W]2f.YY(Z1R
1UHZ_:\aBEEa9;Z7@Q9P:T&?_06G3g7MZAC)MK1_F=1Yg0Qc3@1AWYdNOa]<E7#0
6;2?[NIXTIdO=XF9Ac7-YX9J3EH1>3:O3A^(d.2E+.5<_0@VS5]D_[J0D;N=E(=S
>^4Q<_Ec[8FKcFFNHK#T(#]R8W9gU4-OHH_&N8cSX\JW#(^:P2,7#g:XZ:MW?]@&
Y@/2.FS_4]3CfK#2g>>M_@MQ3E,a^<[e2PQ@?)P,[1W.J9TVcXS9(^g[TX(AX5BB
F5:).?S>1VO/10F0D<dTd_A?8B.PG+I>Ze837#J]XV=QXbC1^7@<<bM;SE5#H@M8
D;2BO(dMc@^7b88[+gd_&DI2)S[2/B?3=#a;5GV7NP>7=/7<FYaNI0?A\4,(f74a
gHCN7aFSNb>L0De#]S&N:MZ_L8ZPLXP69<#P.D2DD0gKQc[c5[HQ<,.8-cWg-KU@
a)2>^W9B:6IQA4=W.F.0,->b@?<(742\)]#&M#U>83NNc6P(-9fda/GZ3f3_VG:A
JAdT]06Q[O?+e(Gg#VYCbba9#Y3AN;.AA?/]]g3R\XA<8#5;VFcdO1?LAI#/9=aV
RO]1=b4BZP#Kc.5F>92:fBF,>8SS&@?3G;Ka?0JK1]O4G/g9,:]db?O1V5KNTc&M
E2<@S<;/(bALe3I09=/-Y.6YfGV<6a(<?#cLV7T#Y5Y06QT00=2]cNWLEM)BL.D1
,ZRBKR#P\CM>Sa.HS[)OAa-#PgA,=3.1Md(..^ZaKW>bFg@WIZSAIRUK;]/36L;:
)<OO\>6aZTEeL8)&KH?beB-XL?[2SdQ5=[5,JVC981=_-H=R>?YT5=fSZL].-Q2F
F>=3V5&DcQW?95BPX?846(]W)Z^ag?J+3,MTO)JMEJ<\X2c-J[5T0c.N-fHF=UNO
a<?6WF;c_WdS,<X[\YR2>W#bc90=M9]QgR770g-GcH65C&eFa&AXTOg+L]/3DLP-
[,PS=JR<<SZ04?O_0V@+B[]W9I77O+DP:SNXF)Z\Z1b=O4XT0)0.d^39.Yg1K@T>
)dW=J.Y/Tcf+HR^ZB-Q[cE>X,_Gga8/X,8_^eS4HbW=3&e/KLGFK#3(,cFDMFebO
0@(H^X,RaP3g@>K?eHfaGX?Q6&9]:/a,0Mc^#T74V)XNQ+19[b/?PeSC<\_0KUEN
66]\3LEMXA;)7W0AV=P2Jf[>b(:MdJSPe1aL47\,RM[+,8Z>]#M5M[-_V=(..G=O
LJS[ZIg-Jg>9Nd>VSOcG1P@D<[Y3K_/,F,&F8YU&9SMc-Y:YNN]J)ON5c+gT:R\O
?[UHN<C[C[\;ERK#43BWVDT5-@NDHbZc]J_2,[96WZ-05\(W92B,SH^)+e2B8G,X
82D>^(g@M,^?BeC10P@\(@-2]?,g2^F-,126-^G_W,ee&6OfJC#,OT6#dQ#^V1^Q
@>7aS\D4^(cT3gAQH&DAOC?;&>DK(9F?_[IN.Vdc]>6>8d(J4N&_BWX\QT17[01U
RK-FeMV(FG[F^cP/X:4I2\BX(H(?7PW&QUAY\Nbd:;dNbJCd#B:N:_&TDX@CK4_0
>T-))Hc,WQ]cSZ?F.9&(XM>Y#PaNbB[J#_E;7G_Ob?G+<2(MD4FVb[K?>\M[3889
0Od&ab9X(:;Dc&_4<VBIYK:LP8?15Y+bQBZ39I\@@4bZN4]3+Re/:U0[_UZN.CDV
def^d:)Db<^-&1Wa-YIS6:8NTVYgC?LT?7NB&W[[HCC@6I1Tc]9O/U27YN4E]QSQ
Y-b-U3N9\><S3)4/VQ7fEF)ZXU/O@\8N<:=RUX5dF@5ZCTW6X7:PP?:&,+=W<ZC8
OGMJRA3fV:MEP(:FEM\5FCJYE#4V5CHZD\JZ<3=G6fG-dFgcbfQN[7ZbNS?6\a3H
7#E;?);SKg05XGR68)&WU^7.:JT>BJ)GUR//QFLK97NC(Q)9=dHcb\[X-gA30.<5
Je3>D9SG^I9].TOENE<eZ-d=J@G&I<@.0E/.I;f[455U#\60-+[>K]BMI/7FC=HL
7f/@QaAK-bH159JfYec[BIXP9.OKFC5\+S0;H=FL6[N+W1)B<d06J,LDFa?Q6UD-
aIGT9<XH1,.V@@FZCJA;]AH4=JK2^<)N+4\;WM6I9<_-\]+=+bRKE,3XEII.-?Q1
AB,+ZZ@#Z5a+W-MJ\FbY?2+RDc-FBV:gXZ2OK)E:f&N2DRP@BFT2#K-/fGB57B.P
DGI&AJDf?<1eL,RIebE9P=/T@gG0Z09d,04[f>-C#BcQ-GE+/LY3W79eWVWMc?]S
#Q6;e=WRGE_K+((6)K8\0f7;H?DbY:[DN+5C2-Za-P>U7.F,g(gTM;/5\LNcV2;4
=JOUTA61DL+/C9EEgTB&^/;?OR#]K&=]+G<A,BKB;LaeLe^9QSf2^I]MV;BeFcVE
<Ca.,R;f/,ScHS805cU-;BM8f:ILUVNGd;&QQ/-aN(B?:B(2HTX/:B,M27BI?,R<
0;GZI04BK\^>Ke2>)cgG<(-Nf+2)fb5Hd<3Tf[DZ)1ZN&<UC45e6\G@JID.?V=5a
CaVNQ_,\(82S331fUYdLLUY=FGW\Zd.gRWVF8ec(BX\+8(J0@YP-9&GVf0@,/Td&
FPD^W(NM/51V2=)#XS,MSQE^gC<.TaZKI=>^SZTg4U54&?@IUX51/OGJf38F_]L5
F?L^4@d#/1+=gLUG[aMg/aT#A=JTZb+ATPGf,OF0+5I^0M<0E,G[e-N[f:M4+A^;
Q/F4#(Y8HCgXB#_4MI;J3SXJe>QLd-F[-=eUJP+[3@3\c?5#+]2I-&UP1?>+BWc_
G@]5U)GeM)T;S3c=TKYX&Y16K9_AdN>P2/7/0T]G>HIK6SS\SX0fJOFXU;.)+[52
)&H>5+6OM=;:]bB>,=OZP?b;bFNPM86VFU\L5-V5F#994_AZ17Z-3YS&2+a\6R,)
LgdN-41?X)5^UP-YN^29,AVc<JY@HKfe=]O[6&(S8L1AO=DbI+3+D_fcVG5MQXFg
E#/V]e3[-W.GJ[;1TP?I41]WY>413/A?325<41ag.T@Y#gg>G_,V5)G+c7()JgRX
(>Ld)LKfd[>:@<5EMOK,NW48:L1b1YPU6LG:g\M=S>f3-f1&4:e5_CWeJ5;Ff;SL
cY,8#+X_0P?1MHO0NZ:H4SEcN7,16RLL;QM7XaT(eZ(,<;4=AA-ILL,;>P/PT0&\
5c(.N;XWUYF-fX;E:\CD0NCJANLeKHT&_L,>:QgE@&S-=_gbQaNUFXBV;]KaOM5T
IcV]^S6BO76]BZRaAg];S04DZ,)Lc<e5d(;FD6C8R91\/P,b5O/IYB&DW;]O/VU)
6,Sg0J)3>e\N;SC7B[9WNLUg@J/IIS-T.)\46e1f[LFAb)-Y86#(<PEfIB;@W<YZ
RSJSQDB2f8Ze8[8LUaNQ8S=Cg([YbB2/G?DS^_4\_df++@1DPY27A#WUN(\#>b>.
OQ?,(,Z;B=cE7J2ADQ(aW4FKA@_0dF>FP.KPS?34BY;QTGZ.X:1,.I=\:--A\,:F
XQa6?_F^ZZQe-G>&Z,gF2+LBOc<#]&#^[R_^0Ld]6)dcYZ51&>XYbJ<^J4H&K?,I
087:aAZZ+=;;L;f#@BH##2:4N2>/HL;dNQ.IeXC32&R9PG@N/_=7XaXbHb)J63R6
S(]LI&T9+&N_0J62Q=L[T9;+H-U>3Q1gTVF+f@(7cWO^&;VD8[UP#Q)HfT,1#aYL
,3A>0LWR/Pf;F5@<?MST5@M;&(d-&U14B/FPbD1,Q2W+,ZJU>deQK7XG(aca>Y[[
]9MWH^&AM6_-BTK92KVMeN>LJIHXWKILg,P8LZWX_TR\,:\YK4^a4D=>(dD0g,17
E1URb<OD7X+IJ16^9D=<IWZ4B35<EdL.37T2]YF<A^[Q.)3J?7,X^c\IR42][Ae4
_;aHa2_cbbEC>JNI<W10S0@9SK5F.=./:5X/^QZK(L6WC,JVIED<HdcY?Z98\G5b
=RK:LT.SUXHS&QNUd7e0]QM;]V+QcHAf&QU)N2TFF_3C\>J_cACgYHNG:=.aA]:6
UAL?@I5?J=5C0DUYKQ(<#cYaFV,:[Q<11A^Z,E5[51L_:a(E\16.@\-/1RLB[)V_
_O[Q3HY+2a3Z?c(dADeb,/ZP2gMC5-O&JT7]:\VU)dB/1a;)_fdd@Nce:?@W&I]C
=g2G7@P7?dU>/\^4;V[[P5<;CbC[-G(5/W3J:<c4FYIQN0VW2L2bRJcEBDO.O;dN
=g=C>PWF=+W_4Z@/F84cC#Y8@R>@RDY9^>Q4A/BU69-R\BF^/a\QQ6-N^b?(-X<W
:b)g1GM(:@7)fE&WBGX_U_T(6(&PKXGJZA#a4^CPS<XaGCb<ZI/@-VbWZ3-/HSJg
S:B@<Ef^bCYMW9D0)I-9\ZEQ=.MT8,6Z;g<Ce#A:Sfe_-0gG0a8f]-Z.a@3f)DJ3
[-D7\IS@X7dKH+SPFa7ZPLA#()N>b[1)?SB7YLE&SC=[ACVI7^Q;d&KBbcY:e=&N
73U6Z(]e5AR/SBO>JQHb3D5KM3G]:.:_//P2JM_6]VZO(d_#N<RbWLFF0S\K>-V1
MR?OYR0M_[77L0DWMK&G_F:;KZTaJCP#Q<EK@>U@./C@N3e@D57D)&S5]NA^L>P2
9^^Mf7DS[1LQFSaKcK(c,PE>FECV-aC<PI0\]e+Y,:A#?H;a4Vge)EgQ#41;D=;C
_Ne^U;T<UL/Q@1AbUU=V)PKd[2OFe92#M+J]73bFN[XA/U^P=fA_aeU1;NL9@PaG
AC>?1QWT1bWQcC\F/QO0aeL,=OFX&N_((2O)b=XFO?N;^dPf-U@2OUXeR8-RVD20
@KM6cCD(+-cK+X^^P6A,0>SSF?He?M2/WH6&1@1)DKPHJH3?eLbS@#aD/PJG0f08
>\LV;+<IBPWC(5,&DA>fb39QA-N;9I1[1WH8V^Y#E[Z0+I]^<A^C9SD;V(JUGCdA
(G,A(g1OK?^N>>:gNXWa[@\;ZD7?3J15gKC(H;71>Q@TdUUT.Xa;0U.4EbJcfU7>
P,^e851+2b6>XRFcS0XVbD72TC;58U61>U&4L0)O]8]-+b#FD)2#QgHc<0Fb3T]A
8S^dQ8?JO0f50U_;+3,S,)I[K3ZYA[-Qg&@_..LdZ_AgbX1(SYZ&ZA5+RFBH#a7/
@cE(J+2+CPNU9_+N#?T5_AbGR5_,E2(XL/bFP;Yc9Y?A==7R>428+3gKN0SLY_:L
#b2)<QDB3S]8NWTP^dZF-?EB1E9GB)RC4(T6J-Pc7L9YQRc-a#.4I)9[#EN^D+0\
d+F5a9U(ZU.f7.#9G1I5<C?[:?M?ZNZ<)K<86?2EJRD4:Z_+NR>DK[]QMWSIg^_>
dZLVfB_TDd25&CNe,@CO_QgPJ6REcPDP[4Tc1f@;cKVfc0I<Z])Y5]/2Q-]N0WcJ
8^6&</c9[/0K6BFNg)0[1<[f;Lg;((c#W1eHE(=QG040@Je:\BHb:^<8CNbeXKK4
IO/\Sb<HU)D<NJSLX2;<=;:ZBC2OWg\SWeTAa;:\NTA,cLD0ZUAGL95(L;V(LJ/(
762E]FEP:9<H_Df\2.VRc&<MJMI5>g\L+<FfN-2OdQ>g>MY#?ZYRO/VF@;BJ=)eX
Z@ZMIW+&7M@:74S<5D06//F-@QT6+8cXO8Z]6.6c2Ig0J6O9Q;4AcF7;=E1LcNWK
U5-:8cXSIH7C3_2=#88\-?WNRQPQ.aF/C_FaIILU\,IL/:,69_3()73&K1F(H\_<
aTW+O53X^4b.OZNNJb\\^CDM)5QAT]50]Cd:H9)]c;S]6^\a7GUV)=7F,46&,R-6
V_)?DS9FDT@TYWHAQUWA:TQ?;]=@g-Q-HRb0Hf[B1RF49Z>0Z(T-F4Ic9=cfd>A0
D?@LY>UA1FTc#1]3N:S[[/DeCGTg=_J([VdJOQ@;c]5a+O,R<BXL/BP]^5Y7ZZQ[
@Y;4O-OOE0A74g]N+^WN3T\;^BLG8Deg&PZFe;Hg<1E(Z_Y;ZEaN[;U,a17aKZK\
(5/f^g>\B+Y4IS1FR0f4UQ[^MM^_2G[&T/WcfKP2DH@fKYP(N]KgMd20]e[MBC\2
/9M(CY6QKUHMg#_7,+UZJRF2W;11cL4VbF;MEO<](]K((dL.c71&78N:P8d?<QfB
3d1/08]#?^[[f]3.R\[J#dHSAETG0C/S.bgOW\X#/2Zg[E1)OW:@ObO,,6G3D5N3
_.?2[BgVP>f5(R(b09133R=dB,.gaT7\83PKN9BIAT\feg0PB,>B5T5XE:<a3I4X
YHRXfELKN<_M_O5PBG<I7Qe&A@O3aJ,\L@M.0cgV#=[HVN,b>DG4S;7,^:?,F5K^
gCD=&&,5Ked0Ia6[CRe&I.7AVU3:,H#9NKH@d7bL,;O[3PbE_g5fF1b?5EFFLQQ1
UL#LZ9#)8K2GgE@bO/2&ZK:N-<eaJ,aE:#LAC=6(?OW3PRNYKYHa0&:GJL;:X&[a
NR0c.--2>#7&J=R+:2&/>9ZJJ+NH)(G&N>+A<8T?c<#:#7/=LUdY2@#SgK=S?R:X
aCQ&@YRR&R[f9(8dCR#@IY1/K0/F7D.A,O\)YAS)IZ^7K96-6.\),,f\I4(4/DB>
H)X[ac/8A#Y?V2d^:PdOS.:D5ObR,K/1-5KH-PZ4(T&>CgPcFW<Z15356UcD?JL(
9UH,H\0-8?B<ff4GB0F56aCPeP>Xd6S,?[4I#AG=8)GbEPCA9COCcI5K2@(1/\;Z
#/?9C>Y&GBg_,XAcKHdQ<C.c,U&_/\Z>e8I),((EULb-d32Ybe5F;HL^AY5_H<c1
Z4XV81g&&ABC:R7>OL0MAD;K;cD#;a/fWCYU+b2NIZ?^0;4-+<,UD&a9-9LB3^8]
8S.E7JdPWCL-g]3VODd#KRU4(Q<GN,N-M9<E<P@V?4P#-;0UDWK6/LVgLL:/^^JT
Ae,6^dgLB1XL,O5KN+PN)7=O^8GUFT)XGUg9/fDf5Q@8\;Bf@AJA4E;[9+5#b=SQ
)cJE4g0F6I.FW6N#5Q<F<]dLZ0_.W8Q76Z.>6BHEV<;_I9DB4D^5WGN:d(X((+;K
ZNVbX<V?#=>N&?,AP;Q@=cRX-?Wb;OB^;8V?T@]9D\7&-P8JO2@a#/Q]/^eW@6FL
715_/Z-.T=H>W\O38R_,P[N5MAc:f3N+1SE[4[#Y1aP+EY(.G<[EB[Y.Y&7V?gHP
+X/H3Q&,IZ?N;SY=>GAQ9OJ8>D3e6cF;.G#RgG,A&a+V<V^)c+>8=ZIFG,^GU+TW
F0_\537@&^<,]aZ^,E.PDBg5HS.<^^Z8C^3G7)FF9C[L.gM;][]78@B8,;/<HYOe
9=Uf,e=)I1S2/6d[G&Q&T,=X(7?G6>c8Z#YVP4VYU1?SOB_7;-U://[\eEXdaB0N
&?Q0UB<@Q.HMY)S2?Z:dPDOY1L_#dZ]>563-GMc+eQ&-&SV/6JWIKMfX@FN+F=7D
:ORdW>5_,RfVFf(HEB(M]NH18BH_<UgJ572fdL[+^WTLE^OX#Id?;R:+\CC:-/OQ
BG?MUG9N871aE]3<W>@RE1-=@6ML7P78RQ,e3[bAed7+=7E3.9PO3@^fVeD+K#BZ
\,<SZG?SVPF0f5_&[2D2/LARFK_#WTeJdbE:44]AF<L?^]aMFRN.HA+fP_?O<BSH
AFVEGBbM]3T&/d5HCF<(VDQU+]+HH44Pa#-ZEA622KVARY7HU@@63dQFFc\=MA:Q
a#fPJ@I>H-<:eP]1e55^@)UL-eF)FZ5YbO(C5CZc,HD11+1MA.gS&Be0/UOc#1?1
@e0OWT):)?A-OYVP-F]/OR:/.3O:LP&V1I@49VTOg#TN8I9?,1S:10dVACGf9P+Z
0,S@LPV.MX]2.Q/Q@O11IEg2BU[a5EE3,B;7O[N\.f.U7R79ga?BCRE0g:L^A2EB
T]V>>a55].(df2)?[1>-#a3C45M+Y;UMKKE^YY2MSc:/H:0dME<L5Y<,GXc?KR:C
6A17aMN]CEJ?1DEDY7_fU2X=M6E./UM<a:=P-fE;\b/K;\HfTTMf&5(LQ3692;?7
<CZ5>\TKT,OIaaA)._R,3Je?-,A5KFU&\8GCUP;[)FJ_&,Y=^PNEZf?[aNUP/5,,
3JSK)/BLLXR^0AM@BDa=TeIX\[6<c.LY;#HU83EK..FC@&-:9,(.+WKTcZ>88A2+
\b5;g.+SCWO]T[Z?2f0D#?c\ZVGH9f;X).RD+Ag#JNM>Z@McN=8/>RV,)/9@5gY+
^Q80KfDf[]SK&/X>=\<=TTO2<QO].?THcDcb(b50:[5c;LY7PQIJ@]@F5>J9.8UI
LUJU;Z(6-Y.a(J<.68SDR,)/1CWfW]3&Y)If,8M?N4&4)VNN=4<&\TN0GOU^;.ZW
XOAJ@OIN7fH<.E&LR2XLO[<TgQdJ/\86:>S0c//OLOGd(SD&<ZR^aZYU2MAb,1A[
R\3Zc@8&S[:;1a3U=ad0FLWcCKfJCeY3I6fQ]D->I8&aeLgd+LOQ:?&::V.g\-3Y
&6]BU@](0K\N2+GO]-X=B?F#,2<aHT7QW]&UUC)H&RgT)RNDgG>Q:0Z0^c:&BOVd
J@5e_[E,P;</f9:7,a)Y1FM(?FCVa[:;)a_)?P0Ba=+2Q\H08e(QUS;fAX)/D+0f
T?I]5.AIFU^2:3>/eOfJR&e-CL@Y4VF_H_SUgU=FCcDJ=CbS7<SFPN80]R0Z&623
fGS[Z5<?.J,)E7C4G)3AARb.X;g.18S-3P]-bDb^6=DY+/GdQaFM9-?0R9<,M1^3
^A>aXFU-K;-CH]A]DV_6TL)g@2edWa,4GO9)E5.F<3TcIg5_V:-;W7BP;M078aYY
=d/^B[55[7aab8_F:ATVE1+F.V.T/=0K,eOOJK7e=7f+X:_HX\eDed2>OJ68_+)M
2S84a+S^+eDf5[GLb&ZRAgEVUa0Nf5.bBL8S3>WPXaRKW]<-7ePLPAFQ&8FM<bA_
:d[Ye_YI:4#7ASR4-/VL4N^?5@eZC]L,eB+TZ;5D.Id/?9Q,V;gb0;g8aWQa&T?1
?YQEU([=&VOE7dRa&FVVT1OWW9L/R71E[?285=R_D8Y,-f>Z,-_B+ZOGBW-;Z.5)
L3Oe@7AMQZ?G59J8??YY&9[1GfTLEeE\a?3g-FDT5&cCY6Wf1XNDYR:X4+:AQ+.:
_c(?X^C0dAg/de--]/=Y:9LLa<67DEF\NE3)(?cVNRaJ2\J&RdfN_=7SbFJGb.IZ
?6@WSM1)Yd_@JeaA3:GG^4,+:3<@BU70]<OBX1EJT8Q1/Q;+L[(,1;d?[+QMSIb7
3JgTO.IA=f;=S,=:EJQD(_XH6(P&a?:7BTe8fgSBb\Y.e\O5?F;CZ6UaNTO8d88;
YKA)+O]031KG8K<[2gWXXWOR2RaU1_[[.BX-RWP7R#H:a5A76&-aRS,.;+cab,O4
ZGEOg@GH#FZ&G,E\bD8IAX4L>,U?]O6[_19(a7J-,2,-g<S:B:TXPdE=UI00Ffd7
U\-=cf7KU[D^<e6)W=3Y,A[RM_c@KDd8YdCUf\;2a6C,Y/;+^LG85[_MGCF<V;D^
Q_:9RF^d/\>fdI>+UW?d44eDP2([+5-^/31cE,+?0ZW.SRT,\c-bN=5>P.FE:45N
]TISJ,_bf]<b0CLeaXRT4MS1_eTSNXE:PRWM>RXPeF-=KPQQ:TM]<;bT+.\SMV@e
WY(?b6Y/>#NK@^EX>B7eU>LGLGK5V)BW<DW[b,7_31=G-T,MELMQ1@YQL^2VEPRV
&L.M-:VQ?O9Q26?]9O4/ITT1/2&R5\=g)XWI@O3VfY/S;THT)e.cECGfe_0_gdOG
7.,C4XQfa8]1U.dYD\\bXB/BMA/RMZ/P+,6c2#:Cg,GK[NU9c8RM;R@JB?dZ,<Y^
L#ZZ/N9I</[DATP@NJ>]/_#_RA7YZ21MVUCZ]a6..LD?MS=GUfS3WHP[1AT1H)+[
g?8TCKK&M-;5\(?-CZ3O[;_C/:gVa6ZFC>cZeg_)Ga,,DPbL5=/aM95OeENTcG+J
4S3H,IE=ES#P<KND>7gZZRE1N[JI8+bB]?Rg>PQ^B-Rf<>0@:cGL63-(XW(0eNc=
\IXb3cJX35OIfX.+RI8H@Kd/2_CJCR;Y8]>M=A,Z<)>1.J.a9.S(I/=6FY?-@]^@
MFd-G(<(SbFfc1(>+>PC@VNgRE>g;O(@8+=9bg7#E7c]4=b&V3E&))/<bK8-TZRI
>EF@5YY,Sd(NTgW\:U\cVa_L/-G&-D;WfKEYGKW7&J?<fA\FJR62_2#G/;aK5DGd
L3fF<-b-8Q:^(d.b2,P5[^1TgMOHA)>@-^?IXb0<6WXC-[=@47YTKH-Va8P3K7T&
?YAf5@LN_BV_be((E)gVa-W.SM?&5bWFG<Q;c@/ba,E69<Pa#X\.S&2gYG#5>TF=
^>0\9ff0-2&AG,HW)J_)A-I6ITCgEY&B=9D?>G:\Hd3a21NTNNZa\BG++QL-d5Y#
]P:2D#9#^3:9TOC&<KPC=P.[Ld0?4.S@=-))9(07G@M0-T;:D)\2dgg(<JCK07KO
7FU)]^E8[#EPdVf\U&PB-FTBQ7BY:^\?BGKMD-Y(\#0B@.V8THP[USTce2e#\5F:
Hfa]->&Z4;5@60GY^O?F:47G5b3/7/Vbd0_+.TI^<M9&3O]0D/^HNZJ(+O<[:@SA
QX(<c9de&c,U&:M6SB+L4)O7P@bbd/b]TeAX:+&8TY>RGCQ)@@((.-_JJaL=P^LX
--JKI(3A(;,b3+2C8B<;#[RBY3(M>e55HAV=HKC_JAb\a9P;TAB)OR6H2]S#/#Bb
3_e3c+cXEMf6IO6c8XQ^ScE418C8=&VEY_TA0U;3\5@-<HAN3RS_NJ4Ub()bBE/-
eT8L,0.#/>2)[dRWCa5?&8K6[[QcCRE@+A2?J_(gJ<Uc,4E-,)cDK/H<S/;OV2S6
^R77]N)S,bX:Z5_992V@RUDD@4B(G2J.GH@BZN9F@0&,NBN)0\+A7>&Qe0CG_f[D
)6&f=;78S3HUHSP:5&1>OU5)U:<C5RAZ3NC\Na41+BN@GFa1)M(D/2)I+Rg^](TA
>7\4Xbe)40M@b-Lf2N+_-?AHe[FT&_W&V6ET(_K>2a:YdTggJ((e?aBaX&[LK71Q
aP(5a0eA1IQfCGA/\7_^:C8>T,7AeJNN4=AW7[VJ<02,-\O5B5F/L&AUEEKN\.Jb
Egg/P,L^OCM-R1&N+9f;^U3J);758YH128Z62ad00UZ&48E;UR618>T]K(41SH^e
E3WDD8RWC,42?0\dCN?;\EfBSDC8AM\I)U9BDgQ;Ba>80RgPS1P4BQ)7[7UF.Tb4
A\@MYH-J#W)HfM[;<H]FVe9MZZ5VZ@//W66CTS9H>[+;7\G;:)H,PBQJT2]-K&.(
#XQ,L=eAZ_OS4U3XW6A,BG=&..EA:D@a=[XJFHBg,^M=T8+K/FPJXe+E\3g67D)c
?N3CZ5^_4014Ea&eN4eFAZM(^KS;T#(;N:)K480)5O+5b8^;6)bbf-\B^_V)N(AW
g^Y=0[Xd2S4f(0)&C<R#6-7ZDL:[RZJ.@6Q0NI>C6>SR4#DPLaH@CFg-.JO;Ncd>
F@BXYYG)A1W5#fb5VY,5QHD.82M)V^8+6ObCcfO^3=_f\;-4NSYF+Dg5D3EC6MMf
gL=R.b.+b/<Td-,b=V:3C89AV>,/]a7?KQfY1&,3SOSS0QJE[Vge45g\O_\SLPQ#
5^6cU.,Pa[VHT\-L,FYaL.N\G7O)W>\H,#6N+ANDIU2I=>=,)42>A/N82G/[@.\b
SdFcO>/:Q^PXZVC9H4gXa?D&O3AF,IBL,R1Q,;b8-ee>I_T4K1Z)IU+L86S1[Ic#
bSHH,6)C:F,5R#bVDLQW_9_4J]@/TLNX)90JPeea#\X_[g@a)G41QMYWNMW?US[[
KOBS&\C[(+J<T_GIDeCVR5XSfGN8V]K)P-GUb?de?AbKb21;K+K80IaN1e3YFJ95
,PZK#aN_.)ST:MU)E0I-Y^\7I+3&4HH(6?gZO@]f/NR(T&Nc:HUb,9LdQR5;H#5+
-)b)R4A5/PES)R0>I\gYITGE7c&4GV0GE,#@bA.Z9<^gg-1.KU8+eZ-9C5KXO2d7
:D6>4B^:K+&(+bf-_?4a(=g]LH]1OGJ/RJ?TW/.I(]\\MX<3J4=TP=<@DF;4[J)L
Y3?#IO?_CI:C.LgM31/.)NbUG-ZSM>V1RfZ^UU3C-UT4^S:@ccI6)2Ic;[cK3__8
Y0-E>I+Q)AM-:]_?=<VZS5QE9LJ&56&0&6T&JWRWcXX7<D8;/)B2^6I<1(HWOZ:@
5GI;N^XXLLCbL-IX/?4[?JORa?Og(10^O<KWE:dNgS]&+WA.Hg6#3a+3EeHRMQA(
K\X3L66NK+g3\HBJ7+W)e[Ga2\./2KYU<WQMgDf&C8Pc\RIgc,daaG61@/R8ZZZ)
e=SRH_abN?]b2/K0Ae3=7bU:A^K:&23&03;,cHKg4FZNf(Y4Z[MH-W2I+429:V4;
V_C4[B^BW0e-VOffI]bO@EBaaWG89B+JXAd+P>DB5-EUQ.IB_-P#7^T?VB=SR669
]:-\_gdP@?a>)YW6_^A(L&EbH;_]:B@:f1I+X7,+0?d(>BFE+KMD-L6G1;P1.dMD
ADg#>N1fS2/V:SY?^3Z<a0dLK;2CE,\f[PgfVV9Z]V/9W?BAS@7a<dcdP8O_<^M5
0g+I;/RYKcX6WeB&+gN)B]AJ0^9OebD>65@[87?4PP\GJ)TD?2bJSK<2YI+967FE
ZF>;e]&&U&[I),-C5KA#Q:9F3#C(2C@Te@6a1WdN][48<e[)&^RR4cPd9X>269-X
7J9^(#B7><B;U9eC/TCRDd9bTIYR]\/aPM0L^WRb?ZUGL^^4Q#GM9b91DO_\5(Z<
8;0EXcPBZHd96_C@<D@QS0g?NAgJMVFR+0&R#O]J(MMM[.A6LK-aT;@.a7]]66a_
/dd79Z9g3/]D:3;];WU>U3c-:RVL+bGOe1R^N6Y5VSb@@0__\cJ3X,2ST\H8g^dK
VUM=.I.=Z3(Y6f@;JD+fC+7A]]gK4&J^b<NHM)DW7edJ-A0.@-Y>LJS_M[WIFF#b
KF;,=Z.RUKB7Q:JT[e1\?AE^3.K,+,_8M6\=@9T#5A<B2/.<DD+c>F:B>-\EDd6(
LM7RRde.N35EV5UY[XA]X(\0>D2&P<9Y+27O=_4VRD/9:PZH#;T-<?&HVX&SUC@V
<_I(Pf5#G_<&N\B#4TaRMHSaAe]5&D>NO6RG\@;^RYGZSf--E#Me:1GYI/Ta)\YM
,@bW5QdNH)/gb-8KWN-^_WPUK&F12SgDU3CI=MF/<H]V&F<f-<4:LSX0HDI?@8=W
=fJW\P^e)+H(#+^,6/:1A+_-7LgKLJHQH3IPdEScZ&e))Q^8gEddacD.6b@<TKL0
MR=<IRe,.&:^^?>#W3PQGfPcfTf4^62,d[MP:9&8?SE2#>]LOV)Z8HMBTOc;L,Ef
V4b6U_:W7g7/W7X/JB:E)OFQ3.Vd:2_b+U/SR^JHYMX)VM_+FWY_BSR=e29<I(Cf
Q>\eI.a5,+Id/M//GWWS<_c7ZN<U34Q,eU[.KC-VE#f]>W1eCEILb\+(H7?[>_#b
-c-S[1^F1B\DS5f2#;aE3.Jg;MRSG(.(>d^PT0NT-/GBJRJVfCf3/a@gX0fE@)D@
Y#_V>3]>68>8:-O9TR\#d7I<DZdePcOHHN2)d=Q#Nb5E5d,A@Q.)(e\1aG&?2QU2
?-Z.ZP4g2/:_@F6;eQSHFST7Y/W(C>Z991B?dAKe6<@eD-2AYgfN00<[aO-#-6d5
KWE;#C##LUXCF_DT59c>.)0?#QB>KfU6,<a6:fUgW_S;eQCP;EI7-MeLSLDgVAfL
XZZ@8E,2RQa?Kgb)7;ZQNBO8HBE?KE\9GUea64=g9;V#8._(^8b0,CU.S7I&/aGX
FUI21PIDQ8MQ>_eO(cDWZ_KBc0^/g(U4eaL>@[USL5,;QKDbVR&B/6AHf-;cTa;2
_MKQOTIW(4FY@KAcX.bR60c/84dPRGa)bHIH7C.GEFHfLO0,[SJV@=Q++dXM97+C
_BC01a\>Q@9]\GVIYWP6YA9I9YL7G_=&T.a3:H8_0J=NMG0NO>2+FYEV8I[Tf#-+
,#L:>\W[O1gV?(g-d.@:)B1I.]9_5_4&&c],I1,_1QI9PLSWZ<XUeMHZIQZSA:Ne
/ea,B&@7TDFKU:eUdNH+/#BRROGZ\g/0Z)L8BS3?gWgc]3SefD:e-?J5)D9VcdSB
BaZ7g5D[_W)M:X;eQ<6b)(8b8T1>cf;<fLRI[XNfI1Z10#E[3e,+@2<?Gb-fGZ4;
&-(TKEP)d,aJf2af4>BESO[)4Pf:^LP76ZSN]DC:K+/QCTMG7N.NSGb=/da&@Z>J
MeTNUI&LC#FAQA\@/GCL:GQ1=+.DX_E_F(JVHc.N.NH:N0VT,d:?M1L)WKHa84I:
X/<Ldg.FR<E(P=c7Y)J4+8P0[))Y_EQ?]P(_[If.V@KPC:;<]LD)5D;-4>(T=4<L
gbM-^1Z>L8egYBBQK3@9];EW\3W4U?Mb0ReF]4Z,]_3LdT9:6V7SB,1HWQHcSCd+
O1b+](801CO\AY8Y9ULKX0d9@/\#;T&@:I-c?_G/7.8ZZ4<DSSFa3E;W+Nc;P5X+
7^-fVLH<c1Q>MdZZQeH.\AO[MdMdU)MQ5.MF/TU[[-W.[UgL9\d?5[[YdKM&QQb<
He;TFACZPF\cPCcdeR7]c;1JQ)1C+)?RZY@RAM</0g8OZRRHE+:)A<I#1S8H7E@L
<R?CT0[=EM1a.9-N<eKXb^[RRF:YT5[^XcPDbCC;XeS;#<ZbAI#eVgb]cU:F&8&E
G,KIR9S0\5&DRJb2c#=&DWE6T2b<TWF1W.EYWg/KeU@0U7Tg:4J07JRN_&^T?eg3
9Na8[?&X])TSADHGRPR275NYb:MA7:/<_C:??W:1P(.FY4R2/892^)>H;84<N:^M
CgF#bc5[b;/)NKW=8JRSEQPD@_f=dLX/;QRHMOJaF>6b4S):fb/AOcI32=?Sb]<,
5F/J1BCXACD7=a&g5,c]2AA#KeU.;2Y3<E,JBf3Td8:(GDTV:SV?b-?#(\XCeWIU
bEB&\78d@-+\]?#e+._J(JR?^)BBE0d=c8BAfW5KO0A]BA,4^(1/Y1EBJN&TH1S1
K^5^Z\7J:NW>Fa\H++8QY;-UM3:(<:dO:/_5+CG@b?HddC&DHIBg5CJT[fDNeL79
:[eT#e@X)R]0UJ^ZK,BF;W-Dd[3cg6B,&;T8=+CQ]#F=ZW,+5?DO5cgXL1H\W75+
N[]cd33A4U7,PL#GA9JHANgEGEaV(+B)#\\8\XKJL[BNKTN9X<U+NK;;@(T:3Z,>
]7#2J525b.9SDa]gRPHAI^(0:TO@dGHUCDR.Y;1U_@6]2HAH&0f8KJN&J+QTR98J
FN@dN:=B,_Eb84fc)c@>]P/;+;L-RHX5H4/SZ(K7J_KSXDfK#.EZJJ;[6T#P4/P6
[)8a/=8)AX3^\^8]a][+JFI&#d;-/I_cGD>Oc_,/]Hea4)_:O^e_9=\K^(X/FeNC
G=I8\V,Dge2>R0-C;09eAFBV(Z.)A#&D]FcgT[ZSNe>5T,Z3.<(8H[QZCA]?)@IZ
\AGcIM9,4CFYE_^^D,0>72SMZ,AHDaDPS3DU9G+8O.K+2eAV@/H:L90-1E(G>N=W
>1UAbbK1=?4f-X3gT#BN..J^UIM@2J#Ag,Y7Pg[-W<VbUaDUA=T@a(b1f6/Vg7\S
1/[XgG\2K@)F;D,aMTPE?PfaI5CH?&+?c^WLIUW]8T=P.SWE2<MSK=O#6Z3./3>G
AS-gd7QOH]VA4P]gN6R1>X#5_XP+NB^&]fH6a5FTCL>S\B>GE6b;M9_30Y>_a[5>
@=E@,VHE)^gR&H4g,ADBPM-HK^9)RT[)+W\Z1=:7J6,C+,_B;ZJ+fe5FMa;^G>@F
B4<d:8A+WC]0bXI=51?XT;KAbZOS=RT=VDaV4JL<39V=?Y=BSGYL[fNa<GH14b&6
2BBZGG2(MZA#7<6JcVQBDAb)F-DR#W,g5(TQ949&,e0cYFFRN[==,.>:)\Q[#OcY
7gF(E-Z<Z)RRe\D<3?GJIY,OgWMbO7M^2-cddW^82R0S7OI>J?A,I&VEL2@Y=?WA
\=NRZ(0FH@5X@?Yf>3Bb^VK77Q+GbZ79&,Hd5>5PF=+]H:=]^5e1\MR]FVEe_)-a
UGL2N<L0U@.S&A8AUb2OfOgg\,-.a;Z+>-)7g(^O2QHV380&)G.WW15RY51[4g:Y
Nb=9BfF0]JfB:&,HO_Q3(#He&HR)dUI]b51EDAL&(a(C2U2ZCNaa&B<05GW<26c:
d?:f1/EG+1E.[;-9[2XZ&V6??56JY8a_WY?;=ND4Td;ND+/d8GZ@;DVK@7R=:BP[
T6<<0;W0=,(0CFO]RU-3RNe36=8N<U^\D#W9T@I:aZe.)@.3)6-/^#O25JD=)J=1
1M=2_([#SPRAQg823XebO]^ML?PbO9_9Y-9=g/2C&VSRDZN+M>38YH&2N80=[MXM
8P#GTDGA3+=ZAP3Na?^?_W5IRZ(]U32-3\_Rd&4>YM9&V__OU9BfM]Z9;/QYC\6I
,AV\a\+);d[FVRdc4NOSQBO0+eI#&Nf08\B9\K^<0Rg(^IPR<QDfTH=LXC5Yb2&7
dHTPWa7=:0\4586:DNB-ge.K<C08PEC@<H<VM)8+g97Q&/M6P[QIbEVH;aW64[]b
dLXg;U4CeRa#7RV/]P0GI&+FZUcIY/_#]PSZ,2KJa/RTB.aEAV&>)&_J#+2Vc=/O
.?P;Hd<-B[<#0>V?)JFaNPPMX^F-J?U@]RX7^GC].LCTY(2JGfH,)BR(-Nc)]5dN
NT4](UW:X7))]O-Z6Zc3c9W:JLC-DFLVJ[(+\LBV[R4ZD8,_Y-\fDG8b9[;>?_Y,
;(?,F:[L@0]&HBV#c[a(#;C_QS\b]Yg:cZePD:(^9NKH>dCI@-XbT,>B0#MEeS\&
:E:]V\M)ZGb8\\WK<7G4=\.5gEEVKRH^.D>@6/f<QIAL&;DfAe?J6=e&68R<HX8P
Ae@:1ABM>JB/X+>NbLeVfR))Z6Q^^^(K#3E#6DBR&5:Qa@STAb_&2g\62+DEU7/7
MaI>>C@C#Y@gS;D;-=8A11Td?>:cZ#9UEH8[&cNLQ0:^ZRFg8eG@2Z+(TCQ].U/P
\dI/K7^:AX(49IG<bP:J]9]B9b#GQ2<RFKFIT[F.<XQ>.3YOD.4_//@D>I)G])_L
B_M6aA66^#9D<7Z^CZ/M-]NPbHP&2=Y\_.?K3I1ER7^0?.b_[95I\9XY)ZN@f]aQ
R38[,5OKX7UH@OZag[b1X#5M^K)42C((1HC<S+R2+4>dBMGYI(0c@7_Q1^_4>#^K
UD?F9^VZ^Y1J.3(]fH_)WK0K\9=^-a\+R:7WPK1,MGW\Q[5J+#MbD/>)H8?K[HcZ
McDg\D=[8,<20N<;IeT/+IW7<:LGQ583XGD[[[9U\#S8FQC=aLYcfU+946JY4H_Y
J:/P&E?fV6N:D2^OM[YWIaF#^gBe+#E7RPA:e<WK2@?Qf;+SIZ>UJ)4NRd2aT;_I
f(BS&OeEge6P87Qg3FI=5S.,7=:R^Cc@,4VEaR=NA3?C9.;2aK]&+EG[27WPF]_2
]Z=O0;gV069NBK-#I:;Of62.LLTAS_b??AeXcO4V;(J(QHc]/dXNf8e:Zb>6Gd3Y
7g>d/L)K>;IN6Dg;AU7gNN+8DZ4,H_R[HEXdcLX@]IT33A5aV/9++HR6eNYNNB>/
HOb&ecK9057@3PafB3KFg<P,KZ:E#CI/6Qa:&FEaX-/=>bef4Ea()YP]fXD7aYVA
9JU8ZE.b.7VUaA(E8H1[E]\:&.cgJ3?C/d,N\89?1<IVLH^U_?O78PO3:&Gc-_,1
\QJPD7IZ06D,\^fC^AIe-e<JDEB/DdX7F2)VDBN\0U;?VFd[S..W<^=>-OXI,D4#
L<GI@fQS5YHMP3F#P\V@+K(O/VAHOW4P]9^5.9PT&BTRAYG=EU7EH#bS?E)>\J]d
ERe#>E;0TCGLf0MV<3ce/YDdaRA,5G@D]Ua7^Td6I@e,YUGG#ZPY8DC<c.(O_gYR
<+]6G^IV0>@gN)V3dE@d9<9S[&]df-ZX=,VPJdaB1<)\f4T\ZQME2?FZM5ZYDX</
7<M:aKL=73b05UI0SVFEgP3gRI0]4Q5B=+WB?bK.0G,F4XPTH;>:DS2J+5\f6:U2
X-P_J3GM46LceEdI/\A<<S\(@J9_8@28/:+c/,R:e.B(#JYB8#F-Pe,ZU7E&3D@Z
?5M;DS&YF.9&IUV(ecf&__=;AU639ECd)FdYYG/:,XVf2:V_^Oeg:?De5,E(.fXT
-ZL&6;?X0E)0:GJg@]bTSLP)[4<bA.G9V6..W^[92^8R<)+WS2H.;02C+2>IY0FW
UVZ]9<_D+I(\L>_3V;=-_OIT3+4(O7)/dHdfRf0Y.c#IK;ge1FOA0NJ8,0)TTY<#
>N=-KeLVR:I^PJ@T3@3Q61@VUS>5C>J#=_WR.:RZN+1>:U2II_2WQ?)5<7LHbBIR
9XM6ZZ\4TDAE70@ZQ4fU(A(S5[^WRCR+..)GdX42d9GO.-IgK/B4F,K5Q.,D>PI)
V&RU1V4=D>TRV:dZECD^41_6@(gHd8C2FCJHHW.C4YdGIbQU]5f6[O;P[689YR4K
4EbeJTRaDL)BPTZd,g;=Ue>3[;9V8/]/@.fY6]XJ_[F[=O&O:/B#5F)11991AT_c
+D:e]Q]6[0;MbP;^@UOIK7_c;aXY7:\B2E9(@fQVc?0DZQ3+C(8YO4_/4&[\d5]-
RG=NY3^7EN(.fdb>Z,#QAgV@E=I3ONM@2=#UfCB]g.]<F):3IX_(Y\_K?(F)99]S
2JNW4G(<S#ATK&-2)aa+bdHSI@V;3.AI?edWN:c,8O_9M]#0cY)8a_;<d((]Xde@
LV3BFcd);OZEI6IR0gKMa(MR]Y3&TIb6)c3ST)0T1)^<AQPT3Mc28:0aJHS2c:#-
c6?bAT,]BFe030Jb+,B4-^Wb@,HH)]dLWL9ObD4,;:/>_/,..2EWPXPS&D0(:OT,
.CUdOL)=DeB,K>0g?,>E&OA9M5=OM8LW-Gg^;.I+A;+M,?QPI\,6_K8b^XR/417M
HDPEMae(N(K?EJT0DQ))]L2?U=KWXA9HE+cKGO9XL(J>7>\WJ0G_dPb96;NIOH09
\WEd9\.^P;4^7b6-F,BI5P6@f8Y_#Q5Vc4HVXZL/QM#JV#1fAAHD2PDI0?#\=B#D
3A\@@STSK[CZggZbQ,&B:A/BP9&C_,X1AaYP3DN-W4^8b.K9a6THP(dOc6WN#PcF
M7NCI-/Te/^<aEYJ;,fKf0/JDJ3@^SDX<WL)?bgBOA^?gD^8JB_G_JWKbYG)B3]A
1f4/K]A):cV1W;bGD6:51&0<=9WS[Y62>2Q+Sc2OYD(D?CY5)#AYd^\:WAdLg(TL
f_H1UNK51OJR?VZe@MFVX?AQ=.AC6#>:WP242GU)K+F+^IU\/eg<0]EUE>)2-61\
ST#=_#B=B)_Z2<.RQ<J)D_+MXPPVa05NMgg0gMgP3,4E/Qd4+D[VH)=#=E,3/EP3
8-3O:>U5S4^a_Eb08AN_b50.a5a;RGYXLE80R0]K_VCcXM882[:1.]FBM_8Z.Id[
24_TU<+Z\ZW9_]/S6QBPOXSTT[U;6WVZ,J;P3dT2[V2H@4;M(->QF-)[T1W&[B-W
ZDWL><8Gf@>bV\L-UO3?NQ:AN_P\6dSAZ9R6;N\]PL0ID._XSLbOA/>0\-L82U]3
QC&FHZ.P.E)H)3?]@=43Yg6?aD0LK]\^eNMQ3XWVJ3/dW=M+9AT8VNe-W@RFA8+N
cgc(=)Y-XJ0V.CL0D\_HXWGYME<cL(Je+T3>1RP6aT_f_d)W^W^@fR(Vef3Jc)S<
O(f/ZYQH_7=cNbKW4-c10a]R[:-?G5\TJUL5=,_]g(IE9QQ2d#HX0AaaI6@BdYDV
CYUM>64&.4=.0-6J\99P>]S01g6O7HDfeXPAda27L=.<OA;Rc,90_G8\aTGZKSKX
&,aW-\fPYVO<6CU#&AZ7]QB@[D84[JI6[N,ZLe,.5REV)??;.VU8LHVg&^H6P[&D
&4IAS1=Ka^dN+IX&LNd?E)gS:W4D]OCb]NV-6?8@H;CX2@_]dCB@D;6HcELVQ9=d
([F?/1f8#,(E#4<E_\O-KKf]Y84[V0(^^]a?M(#[c20CYR(b/-@E]=8H[N.F8U21
eRPY6G/6e1/)-=:Y](AV\+II_b4IYRI<S(Z=PTGEZgXF,KT2MA\_aV6QeJ?Rd;B#
M1MY()P_T2RA)Y.(0g9#0X?[4>C48XdaZSY_14bCcM^?b->ZG\e59/&KLC]f:LWZ
f;A5M=O8fF=J?CbH_G\^\MI@]F&7+4^M)41:]MHA@dC=QI=[3a^YgT9=\YMB:DI\
.UESSSHZ<,=DXY/7#([U9]/g45X];)L>-,B&UKf)188b9c]J,)9,W=eVTaR&OaNM
9@B_a#D]2&AOYF2/#bS0B3FE(T2WH?[A2C<JRB;&\U5PZF/c/)@0FZ(BA7N7I9-\
=GA:_E@L97_NB5a;F(:4A\CUE;<]RcK+QIf#^d@=<GQ=53T3B]6fK/\:GPIIab;Z
249^\YIV</8D]QS^RgWHIeI1+V&,R+(fZ?8FFE:B<W0S07/EQIA<b0S>ST,KMFY&
eH)MW:RId;RaTLe?HXU:b[TSPT)HeF+_W5PNdO?@PR:e]NU5OG\_BF=BJK@P/K:\
+b0E9XUCR8aQVB8D67-NJI/1F&bU<+19D8-[>/=SdT+I+#5f5?QT?@<Ge]e0I;BQ
@\9eX)Q]31CK])?QY)D,#R]DGCag4YG>@5@g3UIQ9G_,f+UUI:6,Jb>EO\fc(Ra.
IVT):^OBUf9&Kf95eQG=9b4)d);;Zbg]>gZfBZ(K+PTS(?WAGMBQN<&ZaJ\=EP&W
dT8\\a&6de@:^cAfI[KYV37R9=S,cHPXe:A5FecQY]-6^eA5IBQ6-f8#f_I\D_GL
6-L/#;XHX?[-#e^-RB^G^F6M_M=W^Y,TgB9.eU:=\,d?_P,Q6Eb^LV=-;6@CVDAS
f7^TQ47R?cAC,&aW&fMfJ)aTC4\8bF>FI=WO#0X,HQ0B]ETRL2XGF@FF;5NGPC4H
9Q(\Z6gPEX>=L^>A1dQ==><acfS-^1a)LJa6fI;>6bd75H75@:MP4\bKB@ER_3PL
7BINHEB^;@[_6<4?_bb&E;\3HTH6,eGMT/#L)[=0e\ROA,-K<==WT1,K0agEMKXY
?(gRT=@>/-La-[PdV&;;D4Z+5PR8;:-E7OTY\)4+#:D2Cf,<G<KfW5\@()#d:G<B
[W,(P/[dJ?#>H<7Z2.#BeUSYYO7D1[[4)=C4cR<,HD5^&:N/P@@\D-JL7ZUPMV.P
R=3<0T:201]JTfJcLUc<F_FDJ2AQ=PO4/]R:R8MPIBWW>c3KM#8WK1U]1[+:fP?T
A2P.b-)bFRZCRKA;B.,G@D];,=QRV:[:Q,G[&-KE>)41&V5,.<Z,V6d2O&&E12T+
]&D0S+f-c[QC.:d,TQe9K[NM3+E<;@X4F[]YBZEDJRN<AQI[UQf#g&1c5E7M48X#
8;b/PDJK[\+S)3,K])A[FBf^NSQ=Y-]]E<UfYO<3>2dT<[\dMIH;1LM2+T@SJL&g
(dEDV/VQI4aD,+aJ>\S32UP(3\bB\)</WL)5WJHSIT2@eT,9LB&08UIJE@=aX+0M
2Ca7J0^c3P)YA0@+BPeESb._)4DMX3OV6DXP,[JYcQ(8.R05:I-:Q+:66VA\P0RP
aMO7Q;Z[>O[&JIdMUa.Od&S]3A<UY3^R?_,#d\,BFD117<[9=C=GSS/^=.,0A[AF
bIcKX0:F/Z.XBceLY].5.Yd.O1)dPNP<,.fY,6@FO##^=Re1O+aC2I[[b15.([MK
1<9@;bJIT).39QZ+-LEKH3b.M77FM[eC/[4IX46/^G\A?X9>U\RQ>MT9LQa\TC-:
&P-V6FXgS=SWO^)]C>>W+&?)9ZVa9e6WdBP,5W\#^cB-GWW?F>+EV@NHKYMSN,^9
<c4WQ._cU,\^?33N,8FQ7OT=E54Dc&gKNg=VV?eP:0AQ/53[0/AU9#1J9X@WbVI]
IOQ6>>Ba2WZH0A&aM<O:\JNf@Rg#07g+7)G<<#ITNN:IE=Q#g>.18,1B3VE(;P+/
4WE])/?(\2Ec.7(8U0AZWM>bVA9WK=4H3.>]/^1Q]+<WHbF]:UD_@=KSO^a^7Z_2
TFKCS?++)^QNWVAW-ROGJR8DbI0E:5a4JgIX,ZEMC;aT<B7\EM+N-#Q?.&KJd2@>
2^a@M(-&8/[[9)Xe7cTJe[3.F/(1eI4<a+Z5,]:c&?:\)UWOPO5;H/<SMPHeUE<C
<FgBI6O9DQ&1.>-Pc?<Fe24gT(@F8L6aC_2&^3#0)cCdKC45G3HGM0B8M^1dM^=+
S>11(A(@<I+)F^>42HO_^BEH:A_[SFA#)C#R)0Tg5e&MKKI15=PX;QF_3E=;dfYE
V6TV&T)-27OTcLEaN6_U_[&X^&\2C[_.Ag8N/D)8?0dDO7@+_\6E;V=)./YGS\DQ
ES?W4W50-f>DL5;EP/,8OCN]E4<38ZBRfPQa<5F?fR<#_+1H1M@bZC@VDTOBgS+Q
^abL-^--2(J:67R?)AfENRQ9)1_H\3Q@N,J:RHKL4P=6JV>6ICG#T,3WZ/cVgW4H
_e.I33STI:eg:BZ]Ua<G7HP1gH/?SDZ2@?&Q&8Sd55AFFdS_EF#3KO).FU7.+]RU
8P5f.1[>&?@-5>c-OT-=0&9a&.D4f>FR<9PYFDAgfS/DQ3I,.F#\U41\9fJ+TT/5
VdC4P\FPa1bKfg4^beK5&<:C6^WTC?KO^dR^.3c4<+G]7LcU:]F(,cf&IL-ZcJ([
13_cT[+)F9/HeWU;D6K6>)8dI(J2)/S(ENQC#^:YKOfL;QbD:SS2):8S8V3=4.WD
P^a+-U_-[b4W<+d5K,8fR#gLW(U74V8LJNb9BAM:6?YVXKTU2R9ZZ6#/)7:53D&^
RZHFa2^@P6;;e<fFWN_EQB:?aSLf(GW&U\^,5f52g/IGSQc)Q);eYJM3>A/0UNMD
,:;e1)]6D-:(Z^6cg,QZgb\T=RF/IaU:,G5Q)S3SYOP@XH_:;34/6:1G6S8?_<N#
&B/(^c9\2Y329M^P#N/Ycf#C18XF9#K8g\R=VLVDIV4E)ZNF^9_=,Ue;=NBN+Z?5
Y9)I@Y1F6Nf1?ULE9[2E]MX1Y\(0.D6Me@(_fX<a;c[KLg^9A.7d>I[_AWY1G\W-
K8YGf6+&B..JQY=U<199AG(Z>Z/6^H=@U640:J#P/5/D+ZGW,YQ#eJ]I?NPZSJ74
R:@ccc\ab)[+0D[JN_KULE8=/=_,GPBL4RYPG]e-VQ;fOMeH[gZdJ&)AR+LC5OdG
R+HDP^1a6g,>-f17c>#BU^JYIIF&V/QH&5F^NH7XD?5KJQMC=7T__DM/WIQ@C54I
J&bT)46:U5A,=9QQ&H?JIa5E][ReT20a[3OMcC[I@W\Z<<D9(<_,KLZW.R9=NM(]
+?Zc?La@;aI&?VYHG/(4YO4-=OaXfLZ&L;L3F[a)A2Nb5GXOe+[O#@,3R2+-:SEQ
/SSK]ZE1gG1&:8a773E=ER:8@Q8^9[e[,gTdU)H9E:eE?>T.\M>7A_Kf[\F1g6]A
Q>(JZ?F,Tc-79L4>cb0e;\/SY2=@H+249&2F]ZO8^A0L,Q/TQOK15T&@:ER7?HVV
4f_LJ;44<T=L-X=#2/^(FMbK^?VTZ5N=@,bK=fH^GI2I7I2MX<0:P6AdUCT14Ub<
)1Q4,(^e0:bSHVHGTA2[(Yf_INZc[GdONKRK-TEJVM@aME@#]HF\W5#=e0KGW)/_
^:=[b<\Z1T(N?4@1G?L4_T24dR,845b[FF#3J[SQU:V0PW^4Oe<(+Ab\@dYW&\,A
b0gf0XP]aIa^a]5aKJ3;b8HT,7^c7#6T[S7Qf/<TF_XD9CL^GVTYR9EIFVYG2;#3
AV<@#aX(Y_V7N-WY))]UBa4eJ19A)NGP#24=M@111fC^H+\W;P6d2;M=XO96cASH
X?e:ARL5WgEI4FH,7)73BXPGdGN.O5Ag7Ic#96T[G9Y/.>d+-03?F&<feVWg<NTK
SIgZZ(3NHMc[/2beR&K+X[-5CgF,gBL9\//@;J&7Q>=a+0(K:daICLHg8G+/9PgK
NUcbPU.V[QE_;d1KYL^RZS@eJ-XSX^&FS-S>^J_@7W9P?T1E7B]LgP:c.JC2H_W_
AC85eX#6#WYJb/X;fW\T)E-]?cPD]D4Y51XC8^.fX0X:FE\GA+W^V9QRZ5V&)G,2
=0&,G@^f^E^gC8TY0-A_Y02eL(AAH4N;2U^a>X2O:]6cVA<B=P&,)E=F2;?2MN&3
C+\+-;HW]SJL.e>)eNM^I@-(NV=G1G16MFD:8#XcADD>EaGY[>GEP77;F6XK2TcV
0]J=]0N><H:R6N\0;5J10.YYHFGcYS/L2PG^HB/g4fNb]cd57YQGZ7dQ@6TJ)V9[
e57GCC4\RD5_0Zc3bG=U5]Zb9VX3J7[].U?BXOI3;cV[YFb#C#KPHf><9@M#+B#,
B&bS)(Hg/36+e-=?HdQ5edFZ[1J>I-T_=-NKK-DM1&c[]6G?T(Y6SLCM>A?W3J-:
DZ]T7D1H9NKa9XOCTg-e_\dbPOZ3dG74<+UJ+8YM.cR^Y8^RYD]ILG?GY>W:4BIQ
R9_5a?<GB>;;0bQNTb;Z&W.2OSFT6C4T<I@[12EGDE6fG;(480E36:=;BH]dVfRg
dD>a<J)KU4;@&4<.8PJbGAST6T)Cb+e\_L<(UPWg\&9L2P4@5^9Fd6fO&1[O@9c.
\#T9>LE@IZ5)LV?,(Oc:Pc3V-ZO8db&65#L<US7&UYd(CIYO+1IWaV0-Y6^G,_:E
921Z=DC;T;9bMg09I[f5ee41S@BZ<;<:@_[-aeAHK>X&C,Yd1DF=cP&(UG>3K:R#
VaePVQ]#6aE&c+1/a-aD,:IVUT:-J37BH4@gUO0Y=Y3N[VN#?ec#267Zc,^<Y0)f
T7IXV#ZFcR)WGAQ(d2+eC#;M6C\:A4PC<#1e2X9/Z;UfU-G;WC.0&AdG3Uc[?YTF
4#1UEK/g)Ff,SIb2YaA6g)0(b>;=U&K\ZdZe?D-a^S_)]C,)U.\D\0,C7\Mc_=_[
5K_VXbP/3e?8FGN=]ef,O[PH_<,aS;B6O=f4?f2ZM_9_G4XOA13HQ)@8&W)b-S9G
XWbQAGETX8?I)-7Rb?G^2dLASG=)]QdKGg.HF=aL&ZbL^,ZP)F?\W6GfI\SHfb[7
8:/Q=&-(ELGECAE?KXT;Z5>N>9R)g>5H1fM1KM\8<2?c?GCU64R0d<CMTF]@;#N1
_+QbTAM7d6N0VcC,,48>1805QYFCObRVcdP>5BV1:>O+<e5@gb</GcKTQ2IJJP>-
_K_1RO0a)=[\\B/>gaPR=Z3Ne[]b\ba9RfLcORS8#eR>P^LD3)YWeeC][5FW522Z
7cdO;H8gaU)Ff:@?82;I0^a?9>8FU\c]??V8;=<0X2\V5VDXHEg^Mfc939L]?5T;
9<#_&V2L0995e1:WFH7+A]Z\V(LgEcD?H-W[TNgD/>gP)>acE=3G51ge4_a<U.:>
9;C<@fSB]INBg]<,X5(CO@50NOQ,SIMH+.E.NK__UGBIE8Q.#:c.PfIB2a(#WX;;
7^8.1P[8LE&J2_TH)2&)H/U13JbJW@^XGL?;>g)M)CDG[daC5^=OX1YW^P0L<Da7
&S+FJ9MLZ>P,\7U>]bU6.bA&cZ3X6X_-G)4/[-1S=BcC1f?,P;QKD_5OGg85=1_N
(&?M\Db9b^(^b>DBA=C<UY_OfNV3Q^9[4S+IX,Z+MZM#X&?K:_?9,K/0#HgTM<0^
JWbHBQZJW,)/ML/OA[AOQ4WAN&^RE^5]Q^N0F0eF;8LD2(U):d+R/(8g2T0a11OK
KG7UQU<29X]b_6edOd;^gDS^^+IT]OKQ\-4\aJR8A5g,\+&GB,KOMRV&KKN7AWVe
GG576+Mb/0@UBJ&>/8IDdJQM5ZTB0@f2JB+eEaJe:H.4B9_JbV32TbG=ZXOD>:4Q
#0:?#<Z>JA)GJ_YR@5^81fKX?e\TD>#^V=Q_bW/\AO[26-[g06(8g4[V;]DF9&^+
-+2?9BI?a9_(J1fW0,YHU85;.@I#dJ-9e^ZO&9GG67)TPO2><9I7IF,-F]JD#V#T
SYNP8/>gC_3=S?\_.K./:D3A1?RE)I+]WeMU@=U,RM?0@<TXST+cKIP_K9=N\/-#
B2V,E;U8&ITP8g-4[;-T6U&_&K>4b9/>C9ba#Od9Wf;GJI,Q9YHM;UU8./G9)8U+
#6Lb.TE3DC;HK&BPRPZdG/9WQX/aGWBB_@9aV/WS8Q/N91_,b@(\c,C+5Z8\9.2<
AC]3fe,]5&_O>BCA#D@[[Q/Ca;ZcPFe<O;F:/^b9^U>aF,GZ#LNI:/+U:/-F\X7Y
821+B2f?J\;C,0B>;AN-^dKQP+]+GS@>(LfDeGa9FfLA),)-fOUS2D]OGCeR)dZ0
&KKHCe]WE/0L^PKD;:I-CGG;,SN3[?)ESbEL@=E(/[P5B8KbQ9(f<9&07e[ZQIe8
/CQda:c;?K\<4A:N:89M#YSPGHGFd+H:=@:f(.0Qb\22W8G8KJdS+0A#HdL_.O=B
+5:[T[a(#ga2<LcM=9N8((Z-LCd-B8g#ZZ?19JX_@PY)N-<KK6K=,.Og:ge\FQH=
MH#W/3]De^O&S4YaAV&##C-YSIG3\=_fO:KGg4]3\]H?dF6A^)ZP..Q#[:-62\0P
1(6:e8a@gSM&7gQ9cD>+Y.@D3Ig^:7I\/>VJKWOML)NY6LD8,C3Y,J3?==>)3EVG
7Y:NbB_Q(P?=H>[X2DBD]aF-S4dSg5S3@:BHIL#XA4>ELMT02;6Z9>CJ3MK-:8O6
7E+_A4))\bd;1X]N]2,L@e/(R1VO-#[E:#-3+2)(,N_##V.)2Q8[K]@[7G.)I]TH
[:gSL<JVV/=01&;F6O1TO61:ZOdM0Q1O<8<JQ3<(NE/,0NgTb&TW=IZ7)BU911eA
?ETL+^[0Y#K6]Q;&Z)&Z><G=W0NBI5V0aV_B5I@gH@_F7ZCe2X[XETNAMCLg3E=L
D701#H2S+A@-CSLKI+Q\#>^\7K&5FUYEeHLNdS/#<(=[K804cT;U&+d]#S5;e=Nd
7@JJUDYUFL\2\XO5#I<VAL\g&3#HT:NQ3C]O-L7S5P7(b)SdVFb5c-F35[-IQ_^9
ZZ_bDf8ZGB,OPd\HJ<Oc)f+SA=V-H7,<eI7GYKR7)2^e7U04X76RNPa5U6;cdZ&&
S,W3GE?d+98NQ&:]12Y@^[Tc]OID<B?c#&H-QfPYdf(:.W_7aUaF\<UL;A(9g^#+
/D5L2a=?AE\O.c0FHafIU9PJf:T00PS?@b,ELYG(GYJ@99(@RZ_Cad_YM21)DBKU
^0_7_)Pg,SV)NZ-d/CaOU3KL#f-SP04?/LO?H+1#=1IOJ>E>:QYg32SQd-7,cFEE
b2>ZS7]+<MbV/@^4daVW@JBCAZg0Q8XNbb39UY,2BEHI8e4[(=G[GcJFES1\)gP8
+?>)VK[KU]TP_U&EZXER0:Yc<Q;T+F:^61664A8,^A2AfI2?)gIE9fM(QLZ>D5J/
cYHLT=I=W.b87A.W,7-fROF8RfFEG>R[=]G16=H:E:[YGX&/3TfU,231G?cKAZPT
6=V\RI>=JCCB-SMUYF8,8AH?b?CH(T:@>RKKfa.DZNW<-E<VO-XU)e#@c=H=,eY6
b]6H><fKM2J@KK(4c<bN9Mb<)5.3-WL+QT(\_;c3GMG9EB#AFA256YOU?JRd)5-S
9=JW(d-2GH5Z8de8Y+BAR:WYd7-NLV33Qg>eJS)^4Ib>f@+d#C5)2CL[1,UD+)8V
V_J3LTL7RN^KS^6-[e7#T#fIEaC=>_WeF0Y28(LaXNMH)RAF7(3.cO0_e,]P;Z6^
L]9OIAB,FNIV^#g:KM6caH9;<L=&V\?Y2-GB#<;7.fd,]Uf]=)FL&fFX.-CA+KEE
JFW:[R-_aP.b_a8NN&E\(<@)[Y4JR#NPa>\eaF/bR[0]?f@JM)e.PV?:Y46-KXT(
-V<-EFgG<bBSYVAI<A9gU;O161fbD9:Na)J[<M8R0A;>2d_V[a^Ve018gJS?I.:T
G&aO[(VM7X/@45^[RAa7gRDB&@+JT5WZ-T?_\>5L,gA8XVb42VU>J8c[>9LdR2PT
CMaX.ZV^8JV<?OcKNQW+A/<gK)Wa87Zb3F0-48JKVf.O,50:2-_AC83[dKCDJP3T
bAD7&#bY+N+3EDOV?Q=;?]+c+7S3I:.>);=^T3HLY-S_cE#CfQL<Ld[^b+80@208
<fC6CYM+++4VOE-=X0:bZ];c,ZSZ2WYW1@aRJ/@37,665&Kbb?c54Oc.-HAN9#F+
-HaYgf#@2\1RDR=6]C0P7A;Q4U^]&>9WgE3CA-+RSR-<=3@CSfA=,E/[g#R(,2:X
EETFCeI;5:(Q])P:,?NZ4NL&062B1aeW;d,/0b#7&c(H0O8CS/R26WU)5&bbK]CV
NBYLFQHHCKJB<6JGR[a]3.BG+9@+gJe=Od;H^EV/JM0R4K?WQ:/.d&LN-KT;G=4c
aMW]d?M6MeAO/BGCU\WRLO3Y_,]N-5O9AI]d.,&2//GK;PGdN/4>Z3]AFd_(Z31\
VPDI:M)W6g1PDJE5==4a+RU2f\2TL\G_2=()842gf&02<J;UO_L6@G)/T21a_I-Y
1M)NW/eS-Z\+Ta;I#0:KS:U\f8=7AN-NI.,=0DXX#<#\<4I8^e8aWS91<HF0[Da>
M4HM&(#-<VXcYORJH(8FdX6_(b6Q_KI&][KS\6U&0b+YFSHKcJ1[a2L8,99c9,fD
?#L7RFPEU.W4JO\H>=e_.=++LOY3f5):GG@fA96YJWN95?_T1B3_2RYGd.-S@UC^
6]]<I47T#g_c86A3N8/4R)5J40QKDLTXL/9]cO;8<AL?LfB8SgeSGVP],dARL&X2
UIJQUI^KTQL<]@+K3BTFHR7[)Z9:YBOW#C=+X[Y:;[.b?)C9R4GP;e5>Y17AB4<X
GRe1KaK+VF.MSCV4D[>0[QEV,:L844FDdI;B1W#2BB@1(MHVeB<^,1Y@/6&T#205
OF#)@6R8]HRVDB4D&IST+>DD;cW4KA7K?-MRW>,af6.,64R=DPUaf=0&Q_Q#gBPB
O;V[H8>=.Ud]R0AD^EAI>OLKFf-,BIGA?LKD:BIL(K4FWA/AG_/aY=D(DNe[]YeY
gF>05aP#30T]EJ\@d6B<FC;<_:&=DOHQ;^K)H]G52=eU&P>=:_U2fMN5@bPZ/=4W
g<eJ3X#(^+:W75ESVc0/Q&g/]P]-LP1;P07+VT&EP);+?#UT)VZ_/:c0[fFP9:;<
Z<=e_N/A#YgfDF.g/@JA2Jcb9e#419<?9)/X&F9Yg.1S(V]QEC&LA:?7OEL[-AJN
OUQ@P#E@X<1Z0-E1TZ<(EQ8DUb>\^6Y9e>5f?T;OYFYIX/.C+=?^gf3Ic9GNRgBZ
7/;UC5CWRWE#7d6\U.4L823[Y6V>+.^2D[WN?fG5gZ4.cKM@bB)Sa7I)LcL=VX:\
#adg1HFAEGC^M;Gb@F.fM@7/LO7>HKF:QRKI0;G)DaM>;&OP/#1&A/OQ8LUa/&=T
X,RT),::U=X1.gHH3^C)GZ:g?QVHHDP_&G_.&(VdD5MdRgT5J0?CdS#5((O()Sf5
+<#HeSV5\5U_,]Z#db:gbD[XP@a;XbH0;3:^U4<I.BT;:]>@E=I?c6BB#M5Z+P>X
Y6EO<?NDKF;>BI8<Y]G,)#6<1c^;cbPUFa#DYK-b\Aa;#UI#BHH8/eT-@:,7P:A>
G.U0WJ,;.cggC@Gg7eO(?Lad_^W]=]-,fU270Z:0Z06]CJCY\D8:SO&<G>=#9-_?
&M0a@G0=e4\+TCDGJ5[L],0Z,(WfB<IBD#=\gYAI(RO1WSNL40&N2#Y#&_g#Z)E>
[2UY,^T.[SMV>+bNb(:e3R5XFO4E<?UP;O.(CQKH]g-<1MO)K,>PGE#f_\8Dg\==
-R8(a3afR6(d>Rb08TP5[TZB2XHJ,d2G=:Hg\KQ-/Q&>DRQTf.@AU&8-SXF-HNUK
/ENeeHd-YZI-?S@>UG]@e]&-__N?PS1JP^G21,CE?a1I,&Cb4ZP2RcTKE:HbMJZX
(:@\6-5M^W6IWNK+3DHMC\F;ZL)?Y;264<YDD3@G]PIf4dS?&^&@_<[)+GSOAO;<
(TFA\7.B\RE]A>.^DZ/BTYcb[WSdK>?K0P:=CbGY>I7.?g(Z_90Yg<004-DPL@).
R<e#B<VX\[bDT<I/aK8GIL,/SD(.Q<=BTCG<^+9DP85UR2-1F5gWCCB(=:BLP/UM
b\\K)S85W@0P]5H>CX[(P:I>&4g=g2UO0-c>g5Kg=6AG/Y5;#0gPG@2B[K0NBCQS
#FX#9YI^_SJBD4DGFZRbI>ZH7B;g<C88L6@X=U5Cg#,S]])NW=#.@&HUHV@?7ccY
3cS56ZCU-1ZUHe]X-b4]=d#cd@RG^QH83HYd,O/F]N_@,eg&3LeI,F>Vgc0QOPNI
40(/KF)ZdQ3[[4a=XDE^9:<^BP_@#I.6c#:XTGT9NM#G[d:01X0,LcFK9P8.004L
BZ;@1\aM6+_2dgB8UO_H(I4GW:-L<=#CR\OXJ]YYE:HB6Cg_dL0:08_C,,KF[(Y,
?]JdNYOe(,#22)0TM:;_78^Ld>YY4G^CWIYGZU0O791<B?NPf]<HZD\83PS1HX+\
/B?\MN@E#=JZ(6[I>-\VAW@HS^G=S0a\d[O5dB#dTIScSA?7U@GU,BT#5Q]=F:ca
Z@aPaEXZ6aS\)CQBL9BR.aACTDD1K9Lg;J<R_KX5I#>Qa)Q+8,B]D-;7?P:LNd/@
K^b\31/A6@@2N3?g0aI[<<0a^9TQX^ZD]8bZ\gC]Q,T[.:GS=R2S;U;Q.,4^)@K?
E.a.-O\45P,N<(H2T7c7GZ>JRU\L.(5SXR5d8EU.U\9FM22c.M^bDAI)R=?K&Z38
gCH2LGga</cP20LegJQ2.XS+J3\VR]U3[((2_X2BbU.WN0/QaIa_7SK4V12>R+DJ
)e4)OKcJ@fDW=GHe\a9?=Y]>LG>OeU<PO&KX&4T#8L/-X-B)^+U1DR/VZ5_A8P1Z
OGRVI2Nc,.I@_,dg=RS/^GLMZ]GOcM(]O3H&WdX6>?\?2PNTG@8\_e?/(+d(N>+f
-O7&S5@bUD1BBG^Q#@J&U4EM=AI5Ue9^&6CaX[XZ_fC=e]J;YPM1M84>PSdSYLP_
_:+9_[U=IF<d7We6Tg/;UV[DB+748eGP3>+7fZYP>7IOW,_Df_YJ.1Z3:D<KC)L7
a\,@1\@[IYg?_ATLRH\5-47NW6d2.S-EZ@/OS(.]bG+T3>.;];YD)).^GaS/\XNH
0:Y[Q#^03U@6==JE#Q4<0O:EI5:Og1g#+WE@:e3)S^IM]#W_]KJgeI8F-&Md,a-6
)W.B&Yba/SM<dg37G:IQ^d/&W_O7<fSYL0IT3gVHIc2@QVQ@YgaK-50;=cbR6SI0
UXZ^@Q3/?/=+aX_Y9=8=C@W3HZ8;L78ccX71?Z)_QH9>?VZ;\>gE64O:-V<6\>O9
ba<-BQ#HPCWF=SDX<CEL^\=73cg16=9\e<Q8.-,3Vc<=.:Tc>]#),-)Y7..B1?RB
2,L]&[?0dd03cE.[)7,#Q+F<1#O6eC@.cS+3^:g6C>:EI#X,6S4.6-/:HWXe]L7)
#g7F;DK1)[dgfY,G?.=?4N54+;&,ba#XJ7(dbG4S/cGg?M7@5ZbNQaNGY><8HX#J
3(B@ed_<82KE=)B[GGX&GR@GU)Ree8#VRXN?.gX1I3(\ECcJIOFC(46Y,JaIPWI+
?]^9O&PMEe4/#@TQ_eV5IR88@+RC\\@_+92f.18?G>g,&<L_@#C8C.C<P<.7WA>c
&^ba<#JB1(JIDeAD(GAe1+c]VQ@^[-?g-O7g.QIDFeY23B[VcTF3RXE#VE#eE&1<
bY,X7faG_-aIA\XJ^)5H8ePKH>=UG?1APKYaf426/NZX^LH.7\+H-K+SH4:.R4PW
4Icc7FEd&5PA[0Z1;2:#U.RB]PP)/D)_+I]39^bXFFUKg-^N#=>-BGCPYCYS0GB8
>VHQ\+A_OSZ>]E[?V02M&U+H\4-G-3GRVX?-=7FXMd8;NR>;LK(HG_2N8MBacF/B
bW_ZM^VWI>3RL9,+2\I/B3N.P&IN]Oe-;;FJ.-=d^BObQ&d>Xf3.E<FCXH+^:&Bb
9HD\WN)SH1Dc>GfYU01#7_L,e.5U@V;#.8D5S9KC::c(AgKM^DdKdW_WZT9G@H#d
#<6FHd(1#GAB>1_6]LbS\>(IV;:(@6Z8T,GUF1UJW7DD:S4T2+f-J\:?CRdDTTc1
\5VA5QYG#W=IeM&EI#_c&7[2M5;BgG73+c<LU]MgS[6G0.Q4OSWa7W^<6-;SUYGH
-^4VGSC\98.2g-4#?A=&?aKEIO6A3Q/>bYJNXR9EEBQdg0e9.Ic(RFTg+>M\Rb1G
;)NZM#+H).c6>NY+@dS&GN-adDUM5OQFLF&IVL)3+TJ;N]RCXcU\5WF(PGA5_.SA
+QF?S/4W[6<A06[)AI2./6e8U8R=7I<06ETR#)L]BbF/0Ld&SZM&d(BP.^0+IGH?
+JR;G@NVd>P[M?O?OMVZ,5D]L.Q\.-GRJEW[UeGcUU7N2;WATU2EA#[f@N&[M8DU
55VB(a(X@aaYg,6f:g:PJ-aZNMX&)gH=R3c8IL5T(R?YBTgOd?9A.>X0&_,g4GDM
2ANa&5aE06/Y()5g+((641,A57V,TLeI/0a7-&>1Be==2cQaR]g8AFbU3:f&<eUW
4^Uf0U<bCa+CDZZWafAcRF3VF6-[1d@P,5;_c]<PW78^8HQE[/cSNQ+cO0/@\B^K
T,A+OUJQfc^7D)3OPZaYJ:_SK\BJ8He=R#Y(>-^9E>[D>V)K[UL1UA2Y?Uf^/PZT
;9UgMRWePB)a7-@)0D;5C\HeJP?HXA.(fHb<#N0Y[G,++F7M7.KL#eY0^?F4:PPS
#@<7,c.F]GNHWJ=XO;d0SW081cXNYFFcBSZ9Y/1=7H_I>=1(DT=-Z/\RQ[M]GSa)
?gD-=3SQS/]\6gM11&=FYL_047aG;eP9R>-eIg@XJTM&W@N2,g8(<c8I;-7_F&<C
&N4;gMeJHQ?:C+J#6(>-J>R89)HM]-361Re5cTDOaIZ5KM=V2bbQ#5BeBg)[_,]F
?X5Ud&06:B[acBa>f2gPO2d2[8dA<@A&RWG^?cSUR3YeE-6BQ(0,T/M+aO:@ST3;
2<)85>G7KU3EE4;c?ND70_(W=KEgU_6a[g9#5(c>7M+a\6^7.TOc72,J_([Z#Rd4
DE#c4#AIM;8EBOB.7QN.g,S^).939Ma_.&4D4Q_I3N@[>03JT=-P9)6JS/54(9#U
dPXU4=Q84R[BT=X+5U5.;);?-Y8\O07ceeJ08BPHFG:V=JR97_dD<],>4O]/]O4g
DX(O/eY0d6^V4P5agdA@J\dCP^2)0J(IRBBFT102^//8f,@Q-SR0Mc12^>#eO&J2
?(A<K9P5QN/V8LL6W@ARBMEJ.d#VC=C(&M3A>#8:1eF9W-cU]Z_#^U[PV?7dY48T
187-K]3f74(@?C2K@@A4WW\/0UfSDLd-PWW5A:4=CN:-QKCHI2^S;GF:3PF/;LO0
^<\[Z@]VYX+0/W4MS1FT?R#fY[Q>Tb&\YU9]IdY4&6^X.:(=N:O9_YBcOC:2;d>G
(b6SO:Y@XHE+E=FYPG98SIcF/gW8+=RAUPQCHD&=SW/>B]B=;eMKPgJYI+/Y8d,W
G<E[#+/\U7a\PC>C41IL_:e7O.]<BC3:^3^L#<P87T([CP.3^gXX7;e]\\/Bg4EX
d-BAYd:OOFd?)CcSPQa(_&.PUc5HK(S)g)NECL#OQ_Fg7ER#7g9VM9eF9,N/_IP.
_^TddMP;,BDgNR(a]=NG_/RL+6XdTQQ=Y+?XU;.0YcL-.;INfWW]cIOe2cc>NJS5
\>V3?g\92L=eM90#H[<SN:\@2#g&#c:e5aDE3YNQ;\3N,:Qd9,#P^.TOV?3>:7d;
6UR(NR;A?^UD6Ug;Q7[4GO_\&D;<aT(8<.8DK]1@+JRB?4@I35MC3Gg#8IN.#0WL
fY5,/b^bcL66@[K&d;069E(WM:K1+Y;?&IX2F:4\VI5[V#7E:Dc7_I[1ad)RXFA.
O3/0:O^cINFX[,;<M2QOHC?Wg;.gE\?9=(g(fMXQ;:<F=BbO>U4(\-4B\#a0bCAD
C_VX_P<a;X\0d?E]LB&#D[?#Ig3c<@KZ>[XU/C?+8\VBO#^8R>)gM7#d@?+HU@[^
A+SN;2gTIH9P5C/=2C]IA;,S7P-P6MTFPWKS?WZ5Of&5.?14Ug?C=Z5U-I7S@(@g
7RFV<Y4?d=T5TLTNE14gLcNNbY(+V9SM:OL)/XZ9O>3<.,&6V98U,TO77X6\KA?,
Xd2MFN\SV1ZIdELDIE8^7;5GGIeU,cP:[WZ[+Z;(IbN]bV\INHB480?IV)C[,8gd
cO=cFVFD1R=.K=RTQ>_ETdNTKLKMI&VS2c0H4(OC:@X7,.V[L.&0=cCbO+@FM:#a
K6<4295R=U)Y0Y+/\04[&M\9@Z\=)FTJE7]]1TR>;QZ3e+FDM3^-+,:f?dDJ4cLX
)^INDGJI<a[aQ?8YL:FNe2P)-42Jg45c,MG8#SO=;#B,a+L@@1aB=JTg/RH&@MI8
d<W(JYgf[YRW,XOdI33\2:fKS/@=B18B&R-]9U]fMYT.WZ=)FJ]SEYJ=:YCa&1OM
PF(Y>9CbA_-78:UD\,:]5OU9G1,)JJ\?QTg^WbOePT)VQD4U]<?M:QO:0+Qg<NgN
)5C+:[,>SC);)C7QYT8-c0?IdYT\L7eWL&KS>SUTL7g)PCUEWN:^K=/.3BX>N0\g
N\IN)RA3gI&7Vb6<N65=B0T3I,T8Dc.g8gFA?PH,Z<VZY&US3BS#WZF8SI>6+RN=
QO-;+-(3^HF<J_)0ZV(GYBI+3Hf[^JAR@SWOY=X1<3JX7598^/\ce>6Y7&eHXcQ]
?7::=GHeN0ZM<9:_ZOHC7WXK;5BS\c?\/eAKOD_W^_#?b=VC@U5EcCE->0bF(/YR
#>R;gd8HC5(7I1+Q1P]<H_F98HPbbD1^PI;\^TH\B]F[)X=d]M>:Y<T]Y(-OOICH
aU?WbOPfdS.AKd_P>B4ESD#+-aP8EPR2?a6]dJY:^,/JAb^>XV][H&9Gd(R/C=aJ
d_VL,P+^?YF\DC@Gc&DbR:&:B[B<T[_6;O[>ALDA=;RHbJ)L>W]^D<6VOXQ-WS)b
bKI=eUad&/FCId>#E1:D8Mf\]<J<9@#fHWQ(_Zf>-@O=_:THeX=J#g8_)ODG(>QH
;Z(A/.0V;]H,=6:L/+=>T&/fM+CQQ05aI;g2+NE1ZTaVB,51?f.CJBe:TKbGc1+A
ODV_4:g#UC61.)N^[QA@16LZ(Y_BY-KfG9?@/Of1GVMN74:++b(W.X0R2bg;N>IX
Mc^WX7/JeP9\Ef9\SE44LWcBK[c#N3W?MQ&U(E?AO<;bZ3bOaDKI#Rg4.bQfHUXZ
3Ve[0>=PRd(:B-HM.86df2<\=>VHG]CSMA@@bJM222AQ.U#?NKQ1e4J7R_+((9O]
^1SLHT8W)T^Efd1^^,@)S&BJN5gN4]2W7LL=BTD9:>J667FPXN?DV=GLHU20?X=5
bGQ.QZQY&b,K3T@)RQFf-\-5M[\);CJ11UMCO(Wf1Z#c\VX9g-0K:1.T-7Aa+&U4
ZCcLZ+feG#EK,2C<NKS;)[0&\E;4O#=DfZ(W=+887YM#7N;9?0<8Y7f-)X/8f^]M
9X\[@gAV<.2<<W8S_>0#G^S;M>PIf\X2TAg)HHbR6[-:WfN,M@0)g#1#BUT^f:1U
aPVgAP?Ma40b@:\H#KVaV-#XH7]5K8aM6P+.9ObSS@,ZM;=.4Fg6PFXcBFYIeZcM
Nf8EOK]b)UbLY_VS2Y[\KTX-6#fA5ff[CTd1)YCFD6E<NHEKOe/6=]gT<@^[R+F-
aX3Y]dJQFQN:)ZCJ1-H[=6eG49\;Be7Z48H:2+)VJ#ZI>&CU6\BD/7_W6gF6]().
Xc+XAF>P8HbcT-VYMeU[<R[PT-VNb-INZe+f+@d&0dK&XX_,EY#I+O]0ff//O,\@
->9;-adOXOR(H3WbD,:9DIP^2#4X?Y;;=V;9H>IVKBX0Ge,G<=S?55HYNYY^1U)]
I/GWbA3<L53(_#U?V9;FRG5G2P-18V^Z#KP\T>6(f6#^0GQE/<ZLH(U:f##JZ^=:
a4;BP)6R#T5#SDR6CVW_2&.+XUc\A=@Fd/+=@^Q2[8f7?94N)d^D<?@fdcbeOO<L
[<G1?D97R1:aRKIe2]B-C.Q0Z_::BgY[CN)RR:;HO&BO.&_ETDBIXVQR-0BTXOED
U+;0d#^JTCb752-RE0;+,96]_c<C(NdOe^8b1dGX3f207X4Y6f7UP92^62_0;P\\
18g.S-6/O7O(Dg>&eOTB10YX:)[[,DDE?IfHLbKG02N<ZONf6:]]Z@O=WER_UTUO
M3E<:,&2+a#d7KfMU4W@+KfE,6A4eJFce[_C=9#)G)9;Kg[D<cCf4#FC.W@??GA<
4ObI7VX2-&-E]+7ROW)M8c@2[)d8?998V+H;&.8&(XKE[6^0,9BI2N0IeWRWba.@
Ff2L#g76&BHBG-35_=?G:B-YFZQ_b,]+0=#^D+PH,OBL3_<9b/ATG@fE5>G6>[?<
#SAb.M:+5a>cdO+QV#UMJ.bL]8]DT8&ZJ(S/:4\V.E;4OXIXHdeCQffWR8:VRbAB
IR1H0T?L[g&aa6;b]Z+G6YQ79gT6GY6M5BKNW8\ae,Ga]]TO]2>WA5N5#bNFA;YX
B8)6=ARO^,PUHbV[Xg=VbZ:)^DJY[>X6g@&G345MIKZQ(\(.Ae0ZL8-X&_,0E3N1
,BA6X,N9#ADA;R0D:<?3EeYZUGHVZ/3fWJ7/+J8Fb4R]fdJ0b&9]RD+H9R7??ID&
(a@2RH#O8FU.N:LdgWMYC-e93>BIKe/8)LI<?BV&CQ[.1D9G=1LB-&\.a#M0/1Eb
#+,0@5/]@Ge==B:HB22gMX,OeA.TE&H+3,5C&dH(&V5F1R?]_6&NdCdM6QC;?TW]
^Ac8RFA#UeG5e<@<RdFW1G^E7CFF)=)983?AD\&SIK6A:T=(^<(KK.Yfb=H.=Y52
K-VG3+Zg,6+#:#X9T/KA_.fUKb_4K/aV,;@XRF14JX?Z(MY?B,^5=>=8T[.0#@cL
SNX<cIdf5AM^:_A5.N(fG7RG-(LYTegXC34c+4@/[G<-/4C<+bUDTBc)>]0.>eY5
,dL##.DJ.RQDO3=H1;PaA1TTRTeNa@[A8&G_ZZ7>0PF?B]JV>4,<[a05<HS24J3)
,HNQWK3e9>g.@a0E&?b9Ka^L(YIf<[Q46GQ_-=?7/-Q#J-)46Q3>=-;G/]?;U>3V
6L<>>GgA7)dN@XA1T9[U/Tb;@+U/Vc/G+fbDD2/ELbc=SGKd1g#Bf3:3E01O[-._
f,TJED.g[Eg:3<K/P0F+d8b<\E(EQb\.bOEM:NfaG7Z5PaZ6#17,c-)\PN-ReL6D
-I<1^RTY8]\2:f1UI++>#C/@#;KCH/S@92bPUXS]B#c,5P#<-=SG2cU\e+\:X=K&
6[1ET66=>UHG_B1J10S,L-EgZdX9Rg>2dC;2KBKa?1SU#\A8-UK5_83V.,aK&d@N
#)K(:Rg-43f=9W(-S\I5Eb:&ZeLVBcITB4S71O0U<(SK]-2g]>VI3S?cE[OGK,IN
eXW)HQ\f/HaL1cd@K76aG#^gPd]RMg+X-DK.KFTg:7K)H2[0=T=#-B9]X(;O[NaK
N8FCFZXQ61Caa?ZYN8D:2Y_]<#R2>>7D9HKde0V56bTJV2[,HTNI)H9_DGDeH8A#
(CGV_GO,;^1?L0B;[]SZ;WBQ#Z91\T,@KCXAc8VD3>F]/@>+Td^./U0]Q;]4b22Z
RB_D=US7DM=0QPZ&2DO9NAZK<./.a_733US4&8+^8.3=CXR#RB7ccLa49<1S\8OF
BT_D5BBVC2G)MH,&W@4eZHYJ0L8NeK32cY0]_QB)#4_2S.6>Yg9Y6Od2J[@fNS0G
[/I)f=QHV)CO2f_Wc_9TQ7:6K@fL,JLL[-XGC4-NUd^f]-94XK<U#=6C)+X[CP_@
G=?Y8A12XdfTL&]TTU_3=22=RJf)OVJFS<K\-ZVS;G5JgOe(-M_cKb?J3Hf2[&fX
WC)Ma6.=aY_S&J--(,SX:;;>g\.RW.,ZP74T:2TSSVe[Y<@[2F=A^\VO&SUO.F,0
2MAH)EX/(b#-\D#I\SQ?N+LQ+<,?-AKLc#UbW>N0bDB8+3Y<EKc^&7a/OcPRV2<[
7g-g?.QeYa\cV9\Q.4(?6=X:ZD&4UdC/&?gP&7\MMG+LA.P7;7YZA)&N=UgdOKDC
f;7ASIDP,KT7S8O@I^HQLUa=Za;)RO/;F@1IF5RCLQX&NR.8)[DF0C_@(;ZBd)4#
HV9+9bV9+bSB@;GFRX7?f,VGW,gYA&7ZZ_L-,@P\bJ3#=I)Q\<5@84Y3\PS#Q+LX
LY,AB[H<K#TTJ&S#)X35cA>?7]3eZFE)_[_I#],YK2Wbd4C)RQa(GH\SPZX1R0^6
6a0HND=8?IQNIbB4I]8,DA##bN.J8&GG<FP6.c+V6]R9&706HWH1Mgad4F]g@B_#
a,g]7WbeB?50K/&df2W@#=842?]d28URTdY(^(8?4K1F9\[UN_O<>]gP+6TCX<F/
O3KR1R3V@XgK_(ZG,D^.MP#045Ue(B0ZH,BDJ.#Ja#b]XJH<WWBO^RFQ/]=Z)(V;
Ge>dbXN-)5WK.-P1#LMd]IdS;W]S_:5,V>H4SW2+M8THX]R=0Ca-Z]bD-J2L[F,#
8\@c+2#H(,a<Z&Q<+Z0WL,b;7cBW7]b=fXXIa#eOSH/<XAd-FBYKbT)8Y9.&TK7W
KNXMPYgd<g3IeA\E\46:7>EXe)c#2RNG?(Xf;?U@>TYC4Q)b&3VP=G\4.,/]Y[<(
0+RE+bX(6F4dVb/Y?&L4;GCB&W=6TERJBf5L/CIe5,;9^YGc@bHY#VK#\O1]LZ>U
A;CT]gI61@R1R#?<W9?.c:dY]1CaX&,K?E4S7?RQ1d1^(9Q0AN6g(1_])]+/=e27
:J/8MC-QXT:F+P@.=2[O:WT#_^O-V7ON5AK<)/FeND;C-#B3ZYO,^^_RaJU(L\d5
SS&Bb,..\KaI>V&)@ITUI;@5M^G[@:C<80+_[e1(_TR?af=0BER74IS244XZ9P^5
Y+P=;^;V,8)\6:MA7Ee(SMVRV_:W)Cgc]0Z8))#Eg/GedN+R1?FN5)B<3IL]]Af:
f+f.@\3g:U<FPZe4[f&>Nb851(b;#]RY(R?=)FZ293\&9#4^422XgM_Q9B</CDgI
MS8YB/ACZD7<15<,EZOW#bP)6NB?\bA0eYDgSc87JJ#fS;Wfg&@_[cc#4(ec53F-
AD1a=Ta_N.\XadZN;4GAM0Qa>S=)8Sf2.&V<:Wd<X>ZM>SEA,/\6^&243f2N@:O,
(#5]GD^7aQZX2HSPKaQ>FK@.N71)EdE[bc[;fcXUN#K)@O)32TVaP_D.XJ\V3P.E
8DNK?b:19^==ZS48QA6fQ9MR>TQL>\JIgTQ)3J,BBRJB\.32/eY.\;g6GEXD4JVF
aPgcYC:RcDBDdC:K&94=T-E#QXN-+J]R.FQ5RL\H4X[>(W-B8>,[6E4?4&3U1<bU
/60ff]cC)9<Qf5:?G,TJfMTe,]6N2;0V#J(+_G(ZbL3(@)O@2RJW]JAB^/]]]:21
4RH+ZU-=eUHcB95;_WcU_:SP3>7<3eRZ:P4HcC)^^>TQI(G\.\Od5WUcMa\[G/>E
,gA1H#J&M@GWTA0Ig4e(G(&3fHSQ^TA:IZ/=e/1>CM)3:5H-,;BGOB3.)+5@#;(W
#[M[]8H@-FB[&OTP^F3RB1:cSG2H@@8RL<C821?6[K[?YS1WGQ35X-d2HGe433DF
+@DeH/VSZAS5##\B/g+,P;C\/A\f:(9(A5B\T&]6I6^/bE?@FKXcd\6=SK(?4?5V
UF>e2V/IRY,P_:19@RB]2RROJ5KX4/_;2V_\M;\U:ZM#IWNS,M)XfKE?NRJ:T>Ia
H(#8VU;\GDA:LHD[?B<TOaT1CX-d&@PB7;ST@L.Z&c5M<8\(N[dVRSM:+/.\MO+D
IH6PcPM=HY#bXfC0gSS5):QOHT&0fQN#;XFU#O+FM+^,I#56P0>+EQF3P4bV(KE-
gC.?+X3GW+K/=gI3NJ?>.EdKPJ)+W82O#G&-;-?<S&7&R-Z>HUI^)IK7&O2:TKbR
e_<@8HDK/E5aKT)JB&g7OUR9S#Mb>D&A8-Z9-C_>_RWZF()2N=^&#/;(:38PG[cg
^&0+Q[I\&^85c5f4HNT7^AF/^;_6LM2\09fZ9,,S&R[acEG^SI@F>/06/)SOJ9Mg
b=a]A#H/@P#d.#MK/cBB?+<c6.e8fX0QZ>UD6bg,UZ4150#PSegVg_=<]3YP9#\^
g0BId_</++dN/<W&0G2Xd4dDf&N+B@2gMe-ZM;H,XOa>QKBQ0Z[S3^YWLb.C2<-;
?R/?CBf858@I3F@daCdc0I91/@K>9PR2S\7P#VR7J_?01_c\=(^2[DN45U@Q(P7<
Vc/T\?WQ&6O<J;::f#?#D6W.AQ45D)cNNK;b#/d#8dg7(fPb)-ObH,@]DU1^3^O?
F0d^A8eb&AR?TU@1OI7=FO5X]/4e^8@-3M9R1O9#_^fJZ(SY9X>.PZ=e>B\-,Pe6
TBSgUI,15MA.)JfYMIH@@R^V[Kd11fB)Z:7=U]\Q4:#cRFNH3B&a1UN3^A:LSGcg
F,33<NZALg/_37;0_2N,aF?Qb[O=[&g=]9(#:YJRK9.63AaZ9VYLV?HV9_N--I;R
,+]3Y2E#GS>,MMfX8;d>NF-\S2=L4g.6=DDWQgTOX^N@L7(f>VPf8L[Z>;H,,VUb
Y.U-..+bW9I\0-XTT<30ZBcYN0=A^:GIH\\;_5B5;NXI_Z(Wd[?[;@9aD4<M<WQZ
+XM-URaR(Q5?IB#e@]]N.UL+O<[^b<W4Y.@eU]?+^7C)8IOK_@1-@fHK;F54?Ca3
E(&aN<ZGUQ@7[4G+IRA@55?b&FgV7G^<5-)5S]fI7Ma.Qd.?PU^,_3[7P&?=HEf7
EN:Dd&UL5J7[H69]N/<D+76M]MLZ+:[&CV/;/_dg_=>M8,[W[BZ-#5c363U<_,]P
VJGX-OWJ5Ce)7+P+S(S(A^>U83B/AX+K23a+?4.S<#);?6[VWQQC\F+P4g,@ATSH
E.W??GKUf89+EE//.:MKe:.WU:8KU=\U:@Za>3:];<Cg_:3I)AR>K[AW;M5_QCfc
YVf.cZW7_NbTP4L]0[Qb?EN]#NKZZ7c;^;E2fA,YS@_3_QPE<JK@##:4[&:;MV,/
?M_6<g@>_:Q;H\);b5(ZMLM.[2-MKOO6X8L75AAaPLVb/fcCeDV6:X8?#.cI4O[K
NFHB(d2(#YAJG;NJ8]e5DYU-A)_39XO]D_4f+&6H;=BF.7?^MZ/@7RSf7N3#L)X(
YPC@.NMW0f>:S8K/TYQDaJ4EFS]_J=^V3_W/\b1;?B&Of^>1MdQA/WDf_Ic3X056
&A,E:4ZI:/1D/\(O;8?-a5IR--JOI6QXNc5DMPYQ.SW1a:fLG1Gf^DN9[12E^3&=
--,f6LdLVTCGAF1Z05.ccX_:9aB<.@S/Z6?<@6J97EfGPPK\_(CIC1XDJ[-Fg32I
MJ++N_U/\IAQg51^YF)()+O]Y-5e<g#^f0DP[=?.Bd,EH8VGMTB-;0/6NJg9#(JB
4V(78DTW@JU12NG6=2:T]MB9bB@-2\4XSd+M[UB]Y1._QOX6=c#E1#g_Z+eR6J<,
>/[V..Y\Q=BcS58aMKbgNB209g>-3RTe?,)UX(QNU-Nc=/UdR&bE9N9=:PRD2L0K
63Ad/)ER4K\.c,=ddOO\3)OR8W[Y6^-<Fa>2IGHD_F+G<]_0/@\,0A8Pf+)G98A9
D].0@Y,Sd,O)Oc5]?Eg)IC<2Z;QbY6NgV(-eNO&?)@:aNXAd)VH[>(DHcU&B?&^5
,c&Ya__>\3W&UKM5dX>Q+KSb>O,.8HP>H&\/JZKXA=M\56?ULG38GO&a[V=RIX,b
PHT,QD-cZ&J@VcO4W?12I&bVI)IYT9>e1QQ?.Z>M9:I_=c(5Y=MU(dJa@D_g?N.@
R:1_8KNL4XBX=-B=-0KX^[]+CB@OY3I(E25fPMcG].C.P>Cb9fX7RQ&)9HA;ROE3
&^=U>,<,dIHK6[5YP#\Y6-AM4B23F@bLR@.@We.EL(dK0KTFd2[>,M5I\F-(E<=[
a]#P&=UEC/E,&\A6MfU.=:Gd\<K&:PM1J#?ODc?IVA/-O4?G/RcPN>SgNIfM(PLc
MI[1RT0V>GX5<QX)LEcSN?gH4G=b837=KT+;/#2,cSAU=XMfF3W9Z87.<H=dQD^?
U2]&J]:T/QWHW#[=c=I<XbS+M^.,TA-2,Y\YegQIb>MSD.]?e,#5&_O5e0:S=62V
C/L1\[WSa;C#,LK<^(RDa]A8eGV8[BeEE,JE@[,T[DKaDHN<>OP9N_]Q8CaNc_4S
g)#<JDg)bH,@8(THN6@B.,R]D0gf(L;E_c=+0\F_>[9MJF&^HP\+D\P+)Se\5=BL
Y\=?VJ20J<&49<WF.,;.MVC?/K)/G]2I1/4<5B^8)9@=(7<7X_1E)H1[daTg7]gC
f&PP>&&:K.:==;0I8#5,(K\d4U;FA?(\325/A7f&D+Bcc1V/I=YIZg]4/C3aBegZ
FQ96BgH53X8<OddDI@Mf(dGg[g)/c\LH9WY5-d;&b:?_#-N.O85PKL?M10/C0eD,
MYLI4DU+GJ1aOF,PR,FW#QC_]\a=-EDAQ]b8#?R^-3=<a^OAG\]NXdXA:cJ#9S[U
+bC8PNDOdU249];-[(8YL2&;+9?TG+2OEOFa(bgN9(JVN]eb>.beZY;a.Y^EKU\E
-g@]H8:_NYX^Hba[_IR@d5Sgf8,L9WMO<RMg,Z=e-3;0BR]WJPC@/H/OP1+\U<-&
SBa-c;-IQ6SU>;XTSI#L]0/@g:O&PYE?\7&[gPGaM>eO936c3Y2A>e0OD?[C3QS#
/IO<gd1f]55;U.&5b5g]UZS96/M3X@T;O/bf_H[,#KNMS5302S_V.VYKU63Q8DL5
Fe);>e.1?ZeS5A[OXG=_8VC9GgQWc<Z+7;X\\M@CgA9JV+Q@,K&)NE7R/XP&/[F.
C44E&BJ/O:f_,4=^=a:YA7+aFS<O3V+UE&8ZB,8?T+7D[)1a3D/&B+e46L-VUH]7
CV-KPS5a@I10NOSbU(.QVddCE8@e:;]<aBVbYXGPU\0_LI:G53TG-FI/_)Sc_1YS
&),:SDV\SZafXA6;e+<:V_NFXT[Xc=B-[3Y.&Sb-:a:O60dRX>3DS&^\[bLT(OMf
JSGVO=a>_DRQD5K_?:#ZD94R;LbMFHWC-2/BC]Hcc4b.;N/)I]8/QXTe1=(;B7#1
g^b=C/B7?PM-.^cgKf8LWKS_K[,FfNB@QDZc.P(R77;Ee&+a:OS+.f3GDR;_6J?>
dS<a/c&J=OTE1#:47T+Y&]GIgLg)6)KFae2S;/M-.Lb^b5,LP^;V;/dJ4KXaC?aL
:Lb@?eO5E4:SIcQQf_9S,(1gXFDfO(+_N_7>6=,XcQeHJ37a<8X[+W:Z4,J4FGB8
;[TJf-X8V)JC[YSA14aE<cY6LAK&Mf23?>3>_7V]KP-TQbSS/2XB.9Ld3GM+fHGF
NGf+^])_J:Xb+QK#&Z-/:G>8N4MNNPf)\M9A,MM(3cFFL-bEFO<b2K^Y+Z1_g9+/
cFYRT4[EeGC.?FQ:L>B#R2PB?Og#_7I-ZVKHAP1C5=g:OB>e4>PJ:C2W\<af3SbH
9-[)6HTf0^dcIHWVET=]\GgHDQ+JHAS6Bc@L@?,2dEC<XIU\R9]&P:^=;(b0YL0R
IUCGF]]>?25Oa/:6OE=e_8?c0?+)c^ZO:Q_aaFG56NC]U8[dD0AaQ^-/L)TBEF9b
9[f7YEcB6WUK=+^Oe1+6PIHP;)&+[U#RE5fcce/Pe?F1HN#GR>XWS-ME@R,LX9f,
UbN+\2S=(=#VE9_3?X4&U\28--]+Rb4&])UU9&FT,37DCJ?S-LAO=:.3_2](cO2_
9f]FZfIFKdM]=ZGL7+DCD#ZB8\@_AK0:>FU6VXXb0eK?.W@1V2a)=06&PU0\5<@N
61&/S^bQOJXZ5UabAJ[EN_M:g/:bH,)a<C)9ag<+VUAUC;E<M&C/9]LaS4,ac9\E
7b3a^HE=e,E].^QH9Z@I8V#]U)0;8SH9[(ES[CJ4J)6(^311DYOJYb.MM9X/_?E3
B:^JF:.L-<T8)];XHB+E]=,-0S-P6FE,W<N4YSAFBbVCABX/9@<.,WMUaDVe4JN1
YGTV9K(KK>6?9RLU<TJdRaDI/W7:&-,H>DMPZ28=78bW/-A:RgUY3/dZC5@J,UZ_
K6A&CDfbe]D?Y0(=CdPe/gO5&8>L5e9P]H5c,#G9#35\gX@aT?V/J8I2G.C_RGDH
+_V).)a2=QXF5dbHdaZBCa6IW\c.K&XG88_=<8AQK,DA[2V1gXd&_=b/3U^g>>Ee
O^L^&M3c6Z8aSO\McT2N=Kg8=O@^Q5=Bgb7V0]@:T/Je5[861fZGO,Y2ZNgY7WYI
<F0;>a_0]:QNc6M;72,\GGFQ\MPM?6b1K8,VPB(H9SN4c;JJ&g1Q5(YRMZE&89.8
M7deTJJ,)C.OWR;B5]B(OH_,cF4N(f0g,c8780fc)I1eaW?,4UL=7eg2/NZ)T)I&
&bL/]JB:HY3]eT+gD7A0Z&+3\U./[L>VBD;;_[6:<#)HXBPb?FX=:XB2CBZ2I0]<
HWF38I?/V=<#d2bVO+.N33CU7RdT^O(\^,-39.J9[PAERP\AEe5DLM>5,>26+fR1
Ab^RCEGG\=_9b@,8)5IP6ZVIcd\N<#M,8;26#dC1/f^-E_gYX]FKH&[B#bD+H^8E
S4690Q3dUE=OA?O1].VEG?B?7[3I@OJ6-MZ29>d<:DAf.aW]ZG7fI0OcMO5M@SK_
C8LRP0a#L[VS;e&g;W+Fc)2a-0XY?&f+V/UBM_1U)Q?MTe2_B@f_GM+?I23XIN6[
U0DB2J[Yc?:.RTVb6=9K:LT&DK#Z^7#Ra_(]FbM.VNK&9ZU_3V[F-U@?_=c:/(a\
?XAZeR]HIKC>3V0L(D.9Db.FAU092P>.__-T#?(<g-LT[?JJ?VZDEN7cTUGGR4.G
d?_3C=@&4Bb6?-)ZD_4I)DN1]:14)#;<JOPVg+I/2-XgO6#-KX;?Q(7VQX,(EU^O
_58+JT6[+;<>.MYgd0LC#0dD#1KH#2+.+H9H3T9aMU,+d_7Qb&L]\?\3@(\WU0,]
RHW,P0W:6N.;]P_\0T9R&]LaL\<,_?N^d#]BLcg5F\fS498\fJbgdaJN_R@EF^G&
#K7Z^?ZJQ@4#<4B6?\];b2D?&)(&VQaY;Gdb3G7BT2I)e&Ac/N))R8OI]Gb#2\B7
c&dFJGOURPH(W:C<_Z/GdZV-)=>:T\P#CZ1.]NA[J6#B((>Zg.ME6/H0]1?RCd#I
g<8abTRMAEF<<E^9VcG]P<:SI<,@3-&?A1/)D+e;Y1:2ETbCW<).<@4YRA:-2#OM
.gE<4g;.?SW0\K.DbTF_0CQIZ-H4#9[BJGIRaK&2cJM9NPcY_<SaeE6S=Z9@+/b-
H;d+dQ+6(M]X-O#T37N(EO>4g0[gK202:IRXUK/8:08IIDD?SD0+FXA<<O@.J0:a
WE>Da=MFPSUfZ7RJC?QR)6&O^VXTRHG7GNH6L9dKU/:gIJQcWEIM74\A3BTbET_d
bK12ONPIE3:42[6B&cHf@74=e;<cH1aNIU<EGCc#-5A+V3Q<6_F?U<8V0NY^gEb&
)9A.65e5b:05fS?CS17]cCQJ6I+Q?e+^[4REID\;HN;=TLMK5\YR>=KHLO(fa2V&
KB&(7E=]8;&?G_68>D;O(TP?a@6F1&BXI/[K4JMg,^=ZOG:D+Cf\^&LcK;687Z2O
d^\a>fTg_9LSd:\Q+4:_>L4b1=HGDD36+AE,^YV;WcE7>OD&cRFbg7AC96=^J(G]
4Z9f&.(g&CCOOc#ZP?=7I=13gFbV8;OfD3_L6ZM^H)MbRT=c@JF<92:V&MI9=_+&
\JDJ^YHc&Fc>^YJ9C@8-<TM?2OP2]=T#.-Bd4-g(-82gBg#5?VfZ+NL0bV99BR7+
gSD9&AHc#QX(,X]Ef.66_gN[PBN:]JTD]X8DcbbA3GC)1+KTP@&:fT.LP4NXR=F4
ISdFSZ#C7@2()GXVc+?OIW##LIa^EOEc(9b2(\KVH]PKD>Y7BU6b3RaC0f7-.7<+
;#A)OFCDU:_IJe6LaU9IAfVS4#>>ZR)S+,K3H_9Db&49K/(<I9.=;8I(KN(a_1:-
QMRa1.e6E&&9BfD29.X7f0&-NcQ+UD)G\UG[N-3:dTZ,P],YCZ+HSE[0&4/bP\LG
Uac.+QMfPb@.\@JcKY8>X?RbF<?/C\?_T^E>,=7,DC&E.440+V8a@Z6.>?#P(^JH
9ZP<dZQ[_20-2\HbP4(?<>/2fL)B7E9:XG]g]4,^[d?bZ^)2)@;ZKD=IUA)\>V;:
;C;VJf3R]YY]V7e>N9U.Z38U+;,+Y_Dc./E?Sd>]X/AEQ:fd:-SFN37O)3=#aH3I
,.GF-H](/b0YdJIM7AG7XR^#bTDJe2L>PBG(MX3DI3:-6W<FSSE-PY/g-95J3[2^
(JLUIH-<U+9R:R^VJ/2+a55H3FeC4g(c[Z\/\EcMQ3T:=:L8N:YV9a)U,UcAK/3:
LXB:P^GO59MEG8EJLPG=FR7:P\D[V#TFNfQ_2ZF/GQDO5(a[Ib)0TW1YY#WcL/L2
UKG#.P-K6B)BA7fde0B(ZC&2YRd)N&e<6dL[R_aff@E9H9Ye[YSLc4PYWV>TV1e,
<\_X2QRJ4Y[?67?MS&.:FZ-^6C?IE^19d5NgI:A)W9S/BN,,[756[7QCCL^2Fac,
/H#CVA52Y6AX83)3A\#8:/d<=ZHgLfCRMNW8?MNVZ7CL2-J&16d7C3?d-Zg4^+L?
4Jd51eGFMT7WZA6EA+>O2f[ARRE-P02fcH0A319R[fZ&FZAB)03S:c44e>O5NU;-
J1cTXZSH#_+A=^eRD/fM\-f9DEC[4RJXaD]C7cRVK2\XbJ&PN-)+=K&5:1\a\4VN
7W75I)?e/]EL]UHPM/fT4OQHQce;Y30A3;Q>R?RP)K.Q<gd.G&RE]K^S:.:eNgTf
C?bSN:(17>&DHZ,D?N3RGV+WIF08=5>dH.S=)=Q,(<eK5K73??_;KV;F_M_V)IO[
>)bANUIY3/e?MT;0Ia)NWCMeNX7Q)eRcLAA//8B0/eX;V3MTG;g/,b-N(QaVf&^R
(Yb/,fb-VQ1;FEETf7\6I8bV/R^(7.+I,T\6S6<cGOPIPZ,HT5#bH0_EW]=IO<NX
J6b5W<83NG0X3#bNKUNH??TRFNM[].>>?TJ&]AGR\g9?3Q&#M686L//DW]:T(A/9
]N[#,Q.#/c\<N[_f9WL#0G#@1&MNe\Yb.W&ed=?gfgf0RM=\7(.)6Hd5b^=-bA0d
2+eSR(1HHO6O@O19c&C5@_Z57BbP:HdOI1e&4c.E@9AG_B>2G07PO.DS=fOBKeTR
&OL/)Rd)+B,NV8R+<dS7]QNDfFL9EbG,/c3a<?)a?(Q2V=V>0650g^+0#+(G20)S
^aQ9I[^@cG>bT4Sb60IVe3DO3E1EY;K7G:\_D_+:H\FO+_IL_8B8gN.4gB._1S._
d?L_0JSIAG\1#W2TZ<NXHPAS[cgW=KbOSbQ>^<X81_5JSSR+bZ946..RAP;],W_]
\XW@QC@F\R:8XIG5^Je+H<?AJ:EP<,_P(MU;\ZeH1gE(SX-b?+gEAS6Ff@)g(1^1
M\aVL//>ZL^]N&SAe#E(8;V0K+g:7@I-,R4\6-W>Q#N_>f,bJY-D.&LPSDb<f;;\
)].Hba>77LfQRJ,X>,?=B]TE@LIRK7^)48d]L#Ye)5G=_]f5,[+7+G>,5>aH])[Z
@dD96OGM.,PHab6@P>>d\/faHL)?JF=LU]HQA/?-Pae05GQ,5</VZJ7NI=eOMVN)
)\<b9K\OVEfQ/764B<[G&&H9^22P,VA5E/2+E?AEZ)#(fYDfQ4>IfJL+7+(Vb]Ee
IP^gTL8X&#W]E;0UaD,A5@K9X,N7?bOBV][_\4?ES6Rd#DdP+]X5^2,L_SY^aNbf
@O-Y2LXX7bYX\Z^CQ5A]A_V8FV4=7G2IbbebG]1NJ9FYb?>)OV0g\g9VM,Te:57X
bP>AJ2b+&P/Z;?HMgBRYf(QLD@ECM#,.IFdKc2#N?.g(5Wg#,.(XF2:D\JgQa<9:
)/.L/QW5?#2IJ5^E<M(#D60&VO@#HQMP=652?4MN(bY\DYNI;F3&[#9^ZB1BC^?Y
_\(e),]bA]&+Y9++],F,NBWTbBfT)YdA+UCA>B:NZb>.](d,&I_\YWR-1Y7L-L2I
.B[1G;CM)S\Xe5+.UYG8V2WFRfFYQBYgP:DBa8IM+L8e<6DbH1J778URg3aC_QR+
SK)bZ;fACOM5PRC:@Kg?WV@J4QTC#ac9(1-ZDUPU>G6+-M\X(3L>@SPALQ<dD/c?
95>O7XU=&1]N4/TW]+a\D[R0OB@.+0SA<VZX1:D2.UOaFA(GVC>EZ+4S8\,6e@_O
7.ZIJCRYTfb=/^4.c.(6T_N@V51JTC6-Ed2H>C&.^85GXU^@+M[eeLAMK6]+16+Z
O^B+H@X:R1FgKND+AZJ\_Z0OCTJ?C(LTe<KD9+(Eb,YTKVV2S;D#LYIHM=Z<KTd0
X?CH]&99E+DSG)V9gN4;SL5\IfT#9[,a-06b(4W=-6\YC4W7+_+f/5[E,5QfRd,_
e0/Y=6]DVI(gI)f#FH_X3(?AKRaCM4X+KdAG:1QNMdFI?3F[)?Wg=):B.WTG+Y_&
A8];_<R7QHS@[YWc@JZdW?7_9ZWHeKYFb18V\8Y(VPC?c^6-e;[d0;EFTaGaYBDH
3F]423=2gaXK4D3Y-56,K&XN&J0CDS:YI<&#XGT10Y_BDCR4(54N4Z5e\LWb[V9I
/I7-Db0]E?WE=7_[]>B8NA.U0KQ=;0UEZD^a4:F#^9cYE)0gN2G,AWd:_7HWVV+1
60.)3-RM:#^^IP3O.T3]cSMJD#TaSZCfGEb\=9b7]+Z9@-V96@B0;44V/QbAA2I_
_cHZfAUQe-VFGZCc:[54QTLLX@1KUcBPb<(f3AHaEL.V2?S\W0-dL]PaN96RbU_9
a)7Ofg@<92)@DY6=52(3dK(=O6-/#Q6F-^g=W1[g+C(g>R0ZS#^I&YM#5FL];1D5
[A4QJ^R76bP@d:e<:3U>^1-1>86&F@,:dS8gRH^/5.2>Q?5U2;TAcRX.eeS5g-X]
/c;9^]DUUO:5=F5bc,DO]FXMG^:HDJ?f&M#WV14@1<b[^D+c3+OG8V1ENd/g302Q
)(d+9a?2)S=&<^__IG/_6>;].Y#)#-]+<fLGOWH7b_=,TSfKPDa:.G0Z>OMG^XcJ
^SNfWV1R,eJ(3)?E,SC0(+<SJ;&cVGcJJT4PA=aF(>1[E2XH7.,VE?++8=,-3Q,a
3>d=-HE>E#Aa[DW-8\R6@S64]^O4K@bTbR8L4+=8^,PaPCD0#Oe<aaM)88RRR></
REJZ#>IYS^L)K<[W3O2HA>H,W?_2N:B@M^#U-@cI+>eJ7U1YN_1R;N@]CR#+4K&-
4,+<D<)W_203\Obg-LU_<[QM,<@b@&CS(CbSV4><Sd),[1/&@B_(:[O]gF43/2#)
1eNd\H7NFZ@+FX;Y25\I>:2S//&SMYTE[:QKBVMS@U3eC@XHR5,dVIe9];-)>LR7
e+GG^ZXgQSU)_H[28EXcGL]PCLI=QD+.S4FfS;=g[;W+579QbE&F?TR8OT=JE,)R
^f?SSI_[;W1YJ1fd/FY,:JKX\K74T4FX(]bB)\dT^-WJeO3T_JXQYfQ=DP.-e#A^
M+5H4IQ(&ZaCQSH,.Z?]BdESa_bUD95X?1XCBGd71(@g\/#d4A5R6F#.7HU+4J:/
.EBI&Md\9\_T<FD+[_+N3W]c;U_2-E&\^EZ<a/>d5P5MR9-E.U2T[-0AaM->eb-<
/b6e;3DGLeB1WHQQU,O#fddCPTBM:KGRB.cV^1Lf4W^@CDP@1JEB:,EDS++2a\\=
J&d[_<7VTdZJQ>/dX8+d\+T<efWN5(2P/L(g-W?c5E\\<c,DR40-76V5?4TKR@ae
#;/c<J^H(Z1.S2B)6EAb:,?[Q_a5TZZW5+U&gDC/=<g41G6Q,?-B(+1gRf)WBR@&
FHVXG2LQ)]>5XB>LRS3a</##Zg/e]a?Kdac11B1+4]=5#I_gT(UUV[-cDS0R,3f1
3+58RZ6UIO=BMN=:IYHcDJ3I4-P=J/6\2#T5K,TDf.eM/+E1:,Y=eS/-SLZ2RaHD
aM,).0(3+I_faRJ)<62LK7[&Y_(7Gf<>aB=?G>+>I(]Z3NKSUG?>bF457ANe<>QR
I@^XMKV0,L+cVI+8eXR_VX[-LCb[71@P&2S&,(eaWV/>5S:=<-Fc0)1=PS[H=EDF
3B7U&E6Rc8gd(3K&T<24c[cR6BX44?=451g35]H(GF(.B/WU/gZ=/8YN;Bg7X#f^
HLC7Y(^f^#1#BX><P<c0G.C>&PF_@GL<,):BT;4^OXE765c<Z4#VV4d^QQgKI\2>
.J,7a99H/;?/@2-XaQ_+IV2BK6a#V2@g/@fLEc8S]L)6fX8?:WIXARZ79K\]-TSF
QL/R1/0I<1cSeRcZ=3SC3<.=eZ8L]AcV3+[]4\+1[Bf1BUPa/.FWeLS0DG]4Y280
(=#X,.CAaN-W[RCC3V1#?1J;>HZQ.5V]V5-F/-JdegZ@PL1<cFSQOAY7?Q<BaXBL
FDL2@A4K42QDZQWC&ZQVR&G88Qa32S4f5=W-bS@QZ855X/)STS(Y\MNBb00.7YP5
S-BQ0S8UIUJF5D-]30;C.:GXgAQOD[B5Q]&;ZH<70XD8#RYT@B[ScNF355bTS4RE
^@Zee-Mb=9d387<L#D_aedZTWY-[B?Q;^(PBf548#Pegg4X04^bHQ::7c-)cL0^J
(M,\&(K:)@D5-I](cf#NOLR2&\(eV2LT98>9IF=^bNTFU>TS36bZJ@0IH=cAMNE/
&BRIBLZ(ULJP11d)Y4],5JI@[,Y?KUTMXc^2fb8_M4/GF4G]<H63-OI<:H^WT&VL
6K?(CB,<]CAd2,/[+B/^NOM7NJaWNN1]KHM6AERUN\S7U7CIO>:-QfKeZ#\UGG1>
bc+-Wa&+Na3_>AE1OJ63:N6:][@;3[/]6BZ5f+g4W6cK=PR6XZTbIZ@S@/R.D6YM
Ze/bd6NfV8[U?@:V]9c<Q;C.Gf&7M+2RGY.HGE1.OT81a@RZI).c68UAV89&KNC5
aN]G0T^1/30_LXHMg,SYJZ@_47Bg^^F3d[^-Zf-4NRKYMeD465fWG4;U\#W9EPKB
d<G@2BK,:\[e#8Q#K-\a4^;D9]H#L,^f0>=@CJ6Q-S1M2PWe2.Lc\aXX)DDS?=C&
9P427:d@LK;5BY65H[_,>N)0(W51&T9f(CD&4aWU,^3GHSCWC7TP?H0YYPD>)0>K
8^@T:eNTE14Q?8STZY:Y_;)da<Y1KL,1+4aY0O9F4[>g5f7bF/(Pg-Oa9&XP.4(B
9MXS1T9F;\=AMK7W)H4La]5HRXAD\K-F+Vg#;21aU\e.8e52=JU1Z=-N39-Zg]SL
33E)S#]^?[#?CR1IPINU+\Ob&IFQ[H4]@FQ2.F78>QePT#b?-AL^=F.5I2)[Da0O
0DJUfEJfR;QS:5ZLE1ROAC#G)>@.+#b5;HO=O]2ZS2>WWC_=&,/Vdd?IHeIce^TL
/abX<P9WGJPJgSZD&=)(C>&7NDE3a]-CNA5TFOYcFO3a7_[(04[NR/BI^b046&25
5a4W68@9F0ScffDe</),J22Vb5&0XZddMbD^B0-SAP>]0f/Z_+)1B2\g1I27;KBa
#=VN16GIB^NWYWb\FIGQWfU0/,EX(A=dea[;9&ES/;?<1M03\0(7.e+/GP36[<1T
^V?3K6f/7IT:-D/H)bD&X<YEaOZd:[HZ]5/#f&X;=X1SXdMX0?,4K2[IX06H@@<c
9/GWEAa\&]O+0f2]2e8fN?-SGFPZNE-cOBcVf2aZR.B4CU5N24@H5R359+fECB;,
O-]#/8T7JD6]5XV+]4V1H@e8GJI5@63^/,C?87AU;H?,PCJG^DDC>X0^KN4ScIKP
)4.]Gc@I4I-0^7<#XJ=cOL1Wa#NKKS.eVT?,N@dAeJ+X_I_^g?8HPCU^(8BZU\WP
8TKLO/1RdOaB;fUSLUe5?e@[Q0(&G.Z+\HI_KVGa-J5+\cT)c#F6eNHd_9N)b_DG
EB5dc1OZ:V0GY80W/LP^SXW6+UQ7M#_=b_49?WQSO#(@ee[]/AJAF6_>F7bB>b,5
[_VB2^=.Xf]O)WLGER7D0[.C9H,#W6Md+F0THV9G.g\+KXYPQD/UWK@DUL6M,U6]
OKM86]<-JIPM\@/NHX0/D5JU)1&EB0<g[4eGN6?MG5F>1LTg>KP:5Q?@&JC>0=9Z
8YK;O6(+::PBR1RSK/8DOREZHa8AK?KYA-VKP8V2c5MV^[6E-2.]0V[8/Ue#RES_
4M:+c^c8>?fa^Na?FZHH-R@A5--W-0YW:]G8d?G)=-K#8C.N7IFd&&-<ZG&S(GWc
Y#&9b\C9CS.-;MAW_-AN86cZ\DM8QO.33QOe0=C;A2B+?fL[#_3#2g69T.Ga>[aL
+QPN#23Se+MSYa0)LGMOTI^+Q6&DcRV_3[-bc=,.b_?FQ=-&BH(JBW^fF:bAb.ZR
GQMC?47&3C4;7Id7eXc8ON:1XDO(ZBP(a#cL(HK=:S&L/3+deaUI6/5R^LC^XWS)
XXe>9QWN5CV\b8M1<]<;4&GbPX\RPWDb8[Y--GGd@S3WOe?(f/JLfN4:&S.VD_:6
eK6cOT6P6S:\N8WX:P2SA0Be1-]EGT3S8eT8Nag8aN)X\\8NRP4TVcA8413).SVg
I._ddb(8LbV\A_JS6V1-TPPL4(--E+9S\WA.\A@;0)/AQg3;ReF50KS94^<D0d?c
VZ7g>&)?:&39(OLF)a#cHVeE)8NXc_H4QN9C\R;INJcJ=T.FMU]<a\O.WKcW<U;,
aOD5ZJ.36f.d25TFc.&@]RG8Nc;-XAIS_HE\SgBgS.>6:egP\+?F\^E;]FLLA]TS
Z)-JN8,BD)SH[)R3O2^NJ#0QLL_,JQM06Mc[[+,=M@)P[8dIgS[UM@0c8E5;a,80
](dA\e_3L7/GDcWe(CS8?9DWOf]-B;AY(4H]KWeP7A;P0TYZ0)Ug+8LK-\?a=5W7
b+>@a[=2YZB\@.WdGMRHYEK?<>VPK3;)b_GN&(>b9eK]_)+?(^#cCN:4Z,0O7L9Y
-Ba3g[bd8Q[K&QV=S^N#6H<:H[Gg3Q8KdL><a:>X]Y2Z_<#eMD_GT;IaC(DNaCVB
A@-]_7We6>gKY;MgZ?NfNP,S^?a;6[_HeCHKSK,7X)e6LWG[g]S2fB(.=MeJ;R+)
;;Ra(M@IWQPO;,FU<PgM:@0Fc9T_I?_Cc^A?O6PLYVSggH&9YC^5Yf03+Y:W@?EJ
GEW]NcCG2I863)_>#+cHROZ9-<_)F\67IHOY93R&/G@KO?OePEgYL3dN@MZEGc6:
N(.HG2/7/BDD01e@fYQSX5[BdLL=KAdcd1^ICU]AbL___M)&@MYXe>M^=8UFfYSQ
C+=@bI]0c&RB)-CCV3^KbXE+P7?;Lf8DXD55MB^&W\-5/#,4.c[>X#a-IfWaW(;J
77A3/J(4GNQd?Jd5->g(ZSPE=20A5e4<=Y(H]]99.(HQPPW:@cZ24.gG4C&\3gZ2
96&JQ/&a0OXZ&7>=4BOMH/5FDWK((Bd0Lbb=NgU)f@g1@;?JLDb20<8D.&=?;7eH
Y<&KVZ2\MaIa7/+[<J]P_?A0IOG=/9]]NO/\2;g)X]PW&)aG1]9bKC#O<,<<7]/&
_MZaf1F8WF+9YUF3\<RM_5AEARZfAf@P>@WM,W+g?1BeUY=E[&JgeE+E@)R\#ZKI
4\/S--ZGD5W._Q@=)K6@<5@H@MM6acVgOUXO7X:4\HL/:=C6aZPY1R42DXPOWXDg
13Y]>I>HP<:0)P&JAQM@<4.-;VYQ>OGK9I__V?Cd:;=fY?WGIG]<2J+eU^>=9[Ya
Ga[ET)2#+E.@BbeG[M>d;W0,a=G5(B@TAIN[[:]MT^N+DD(XX?^O[#JXJ,Gdd0\G
b,&ZYAV5N&:6MFN9Q21C20fO&HI0A[gOcB[=T7LJYW)5N&Ee\EA3]_DQ^Eg]_;Xa
616U3/5;_XTZP9e_^cMDP7f:>Sd[</HV=DRHHaf:(9;=/DQ4.SAHc4Yg<8b7/G_?
c6^3OUdV[-3M&NT6IPY7AI=Z>P152546U/1fO4[8/RU-\R>AWWVMabOf#>c#UKHP
HWL.1[A:8PJEZD<3,I4b+.P;1CMc\[A>^7)@6f2ARADYEU868;W@(G#IT&a)GJ@9
aPY-N[XEAO@:8EQ_a9.+&R88QUNH0/,V]VWE-MB5VYH)LIDe9=3e6fO,_:[1#,2;
URaf-/g^4+dT,91R^.,fC+0L^Fd#[]A;GF7G_OHfR9-A/>YfDOcDdEAT=SW)gVNS
K-,.VGKa\@Y/TaafHL:.<]\3FO^e7EDe,L8E.2.XW;2+#Nc.A0U?EXg=@K(?X::_
@Y1/(HCBgL7YPOW]\gT>6]6b04G+WS8#ZcFa9aQPRP6>gVaEE)]8R#-+PcC/_A/O
LXb:-B8KK24WCGdbe>a68Y_TQ2b]aCORJeLHYd^U,IJE\5Xd5H4c^?\2NI1\D73+
H-I/\^)Ea##3Y>:G=VdbV71/W[I&J,K=:S5N7<,e:8\6;aP&#(KDJLY#MBE[@0_T
U/=3]S4QA.=U-:.YU,Y@2NdRK0[5Y0bMXRP:-F[3PORHagV;8eCgNe[77Q;_eQJc
VGX?5]R57S?>CU4Q_HHBeaVWdR\S7Xc9dCcTJ12YV6^PCd^4O,N3,)C.I+W\,4:]
;0/<.?^YBX#83.8E]FPPTK^BLC/1M?T;U1:+(=,><0GIW@#,^/0U,=_B<5VfMGNe
>&JcKP:YG7@^.=W<=0-(T&4\&#JQ\@b]7>;#WLA5W^BWLU4a10.;.2)=]D[1d0N<
^//\Hg^8#3)W^Q2]I7L\KfeMCQI_f]^M07L]<5#7Z&C7SZ>c>4OJD.47Z:>AC#Rg
9TNfTI=3cYF@aL;8H^\Aee)@cbD#Tf?NCA(YQ1CR=^7,75S)T,Pc8^dMC]8:fOL=
^/Y7ER3:+;=NM8]L(/_?SdE_0X?JK,L/V8[MDO90d]LCR]=MaE)dIeCR@[7J-IW@
b3[WL4L0CS:D(CRY<b[Q;@]0L>>K:7V[>1a\7]JOL^ZZga)YVaJIb(EAS(QP-T3c
QL:W7c08Z=A@M1\\]?(d85ZOL0(f4B1VGWWL68/3B5?=SQc&([R#e-UPVQJ9VA@\
<+<\>Z_Z:?-Y<_3S)@R.#)bD5;WD0D2SL1,=3dd^2U[27/A4G;5ZW<[9]\LVV,3R
3@G]CRVQ(U;)&[>-cFI[O^2Uc)Z<5Z;COOF04?O@.dY?-,1JgdefJBC54feGIBY4
a02(Ggf5C7;\MK4f7L:6f1+@UAK@OL\H]3)PaVgb:8HN<^9V-T.<2cA=L7/TQE?H
KI+[3FMP4V3=U=:gJ(Z26\=UeB,:4B6IcKS\0EQZ6X(.62V\9\H@c?gdC0da/#QY
VDgUJ3\KgDP>/>;1OS##7AUd<a71a\\+J;S&,OD=X5SO^f0@/\(;-##LIC:7J,V9
dfIH6(J/cIQHX45+[^2G\G64/30^/&2RAD07VNQ]?WgZTcbagMSJ08GM[a2?TXOL
IBb[7(R/7XCd:_^,>KL&,C9=)0.e7QFN-0RT(EW_6>N\_L2IK^_S?=@E=RHA9P;a
BT2N],PS?]>g+&5cQYaO(@b&&2MK0G<GVgE)3&DMD:13eE[He+(J(6SegSYCaMW#
97S]#/DD^M3.P.8R^U81-?#DQD<C.YC\A@EcRIP;C&AM<3PH,R)(J#bEP>[3a9OS
cI0_]2G1aUMfEUS+[<Q+9Jc_=7#5GGD0OaANFL@T9B_AbF96J:A?\;=DQ[D7XfL=
ENALR5G,24^8EYPSRd2B=<1RXaS@/CJK79<GBTKcW[V1JV5d=f@CY:_8)d>BAU6>
>>9Y>&1\LMZ<g.&Ne?a[8<&BMgD>W1?)<@<T69PLBR?MA;/O4^8HT@AANZUN[.O)
fU,LO,0NQ0AINCB.K.T;6O-<-O\(O4^6B)Y)#@eLWWTP:-c,FXP3R.H8(,##7#]f
KSGDa.9U&?-Y>TTV&W=6dgEAU:\S/d1gefB/Le)Ec4^f^-fe@@U<P[<@L@MC342T
;898NDS[^cg7&dC=TZ[=g3I_>c_4g.A7+/Pd,26(dZ@AI09^H7V1C=cDH42dfW>>
2.2(M50eYePRePadH3J<\U1HDRV-#5Y#+P.YP5:6d(V];7eBU;c-.X.9E6P.D(10
HY8F+BcKg])?f[K?D76/\6\gIB,8f_Z,F38_Rc.Z&8GA/0RcA^[fZg&F3gKaY1:.
-c0ER1T(dc=E+V<8?0KSW7TSaPY/Z8D]WA:Jg>/QQ^)#/7Nd_gMaW8@/N>\<,UNX
;Xff,G_1T64eUIRc:Ib22fR[]1<<7X6IfeM4H1[gZV>LXY_PV86[#5J,g^PfL;.U
86dQAEO5;+=CV]YcU)4SSEV<?SK.2OGSO42+M^=MOQaP,G-1#2,M1d70(5Q::F<[
GScWc.0RH@IaD4JaR?8bG.9U](cecUJ95;Wg1ZJ:.@G:S<HEfC)T:NHLBKGT>a&g
=,#I?<WD3G/KBcD?4K2V8[A?QQB0&:6_+M>6/06LdQgDe:TUUg5M,632)dTI.?8D
<Te7YTGAQIL_H.U3\,U4B2[^AC6?5S97,&c@fD)5W?WUJ@PC3cL@<26T(&LN>@19
8SALTK^@Y38[A6bA+[EQc[B0_QQ8_+R_dXLSR+]abA<6#P9&>MX&X;<BJcS]AODC
#I3,4T,B8P?RI<cGAWD_R[XI#?=D-KSF\95RYJA(,_IUXg<d.AMTUGd.@cY:F0ef
#AX+>Q\/OK(cR4V,VCJeLWe[=@;?NOE_=F4cPU(D@dfMSD+]3>6;c=/1Wg]@CINf
HcSJXODY[CP6]8=#Q/?B)A+,^S@M1U_7D82c6Q^TBf-,gWdAYdMb56W=A765LM7U
9U[[OVSDR5SM2.E:Af,9<3_;a/WY-40>@T&O9c9)8^OK??#KRIYI77#/Tg?RgIg<
b2=MSLfWG6=J<TJ?G@)]HREEA84c\]F\de_7TQV-e&Q59C(a7V2U<Gf-#Ug&MFKU
ZYBU8I0fY^:@X#V.89;g1<Xd9bO)5;WQQFA:HNG7QV(ZD#8#64;;LELF9LCd7)Xf
6^,DTDB+:d^F3L4+BeR]=I137F6KQYP@(LH\#85>3d-#V2S3O_@VdgFaW:WE)W>L
<]WBHZ/PUF-L<<2^\D?(5>I1/NE8N\]a95[91,3.3B9PPKOPCONR11)W&]f6,4b+
R.8fT&+V<1S<YTC-PZF94DbAb/ZIFZAI._fWAfQ;5_5D<FT=>@Z8d^S_gR:MVH_d
0-0C1-Y:<==+9,\?I53B(.HR^H]C]@BPE5RYEKC>[Wa\-R?cLa,XY1Ka+YFPe-.a
XfZUY>@KE<9^Dd6G3.CM.S9^SA\95NO\U2M]1+4Ya=D?5/9UJ+Xge@M2.8>9c(Lg
XR_K[?UNNICN+YX&\SM6eI(XF&/aZ+](_dE982_16WdS/g/^MRZ4^D-+7@Ke\+O\
>]-(^((Md3_YbQ@g08].9H?:cUed1I@B(4:9=:CXcM9J4(K0?dJba,D0>O>X4F_O
e\bKf(DLS/ga/c/U6W8_WSPW#R^fD9F@3D:B^VYB#^[\E9\B(K],KFAKF<J2;Z#0
M#f>VR>(3GeJ-JRb@UC=:f-8T2_(_g.:I^X=V/-UMg_@(Lb>EZ9Mgc\1IG+.B6@\
DO,83688WY+KN,9HX\0a).?YKGNI>&Y6OS?LcH^M2=>Ge])YGEF@aeAZ9dF+JV;[
9MD^AV\HfRY=fU=?I?,f?\FSg/W9ETY/deIK2S4INI()C_NOA@3JCG#@4WgcHd6Y
>f\Pd56+d?c8)8CZAZaYVKcXNW0Of#\IXF=NZ<\N]HXG]+O;Z3^[:P^,I:X)U;Eg
b54\Ea+.YS2H^UM9/BGM97ZX7X,aB-,?USg0bMEZA?&M,,,P9\Z:R;@=.KgY6\1a
)FeH6&Q3dQJG;^N7F[[K]<BF3>.S?H-]bFQc:2,Oa^M]VAEES_<;]/-@3dA3([53
:3Y@?ZB.QBK&cM)C>4Xea<A.Tfcg>.&=_3M+J6W>)@K>&Z#D9)<\3O]=])I9,f:6
Dg#X)7>aENX2eVSN?#3_W2A\+AP?8g;d_SH11FP.9C3]NSRU8N_DR3K<0]J]3^Q,
@67-3aAB&LXW]^[E0(SO&F]QJf+A-@S>D2Gg_(X0?)^G9^B?<K?@(UBE]9cgDNLZ
FNYE(>2:Q>@5;07SUCEYUMVNP1&M]Q=2:Q9aZI4cYdJ]:+&REGPOR2MM^ZKAB]@\
AYf1Q/U80dJ+efVA@4I<ZA3_]EadNRKGSVHWD7\_5^K:^):IG2PS+-ZLPI-_0TbR
5ZE?IQJ:UgN?D)Ue=cFVC0T1cPPTDd)2;;Zc8>14aIK8e:@?G;U0L&@1KMRP_]A=
HYQ,Pb79Z)E^gG?IB@N_MYO?E9&HHP@X\Q2QC0f:0NIXa^-,cY(_8O/0a@+RS@Fg
gFPI&114Lc-aKT6_=4A.O.H&P^0@PR(KZXZC;aF0eD&4Uf11Qd]:1/+XFbO=T24^
1==\#@aX>]YZ#U:8_A:CbR/5]8.63)>MG/^_,e)/N1?VQF>BMF?b(BPAgdQU#d=.
A>339Jf8HKAUT7AJ)S]>bWA1=CGX/6dL<TJA>3:G)5,YSgFUQ:V\,]<B#HDS[aNf
^8[^KJ8LC<L:__/WaC@f@4B2)R5.C2T_b)PR?P7\(DOA(M3Ae.d=O:F]HFHQ:SaE
L1VCC>C6_;67;36P)1=5(--LTM^EA6\eL]N^5K<KJ\GH:_,I>,XZ^7SLUR-AP5RD
\,ILO^fcK1^HL5Q&<:77MQI^DWd6VUBcgTHFA6MQf:?M_]N&Sf5E1c16I7[&5\MH
[/Pg(cEHa:U<-aK]\G\JLG9I,WN[./2/H]_Q.VRcNc;9:b_YD\b=MTR?95N,F8d/
Hb/9;bS0[[,.^B.R[K)6\9APK&N3_7#Re7._9V^Q05#6;/;6RA_@;I1^KfU#VVL^
>0E4JWF4NMc4<SH^cYQWcZ,:1I.DgTDX&-?-#[FSd)ZG@e]?<,67I;Ue,aTPKbP8
4.N\U6c#,2:=@(EB;LDMX.e8\c,L5P:-3;50RTK?6Tb2\#>L]XdQ\#QSVe8^^0)Y
&7[S1O=<V:+QK6=#+2K5G<N:^PLD6I?c[5@.fLW(>Ug<+6aJ3J&T;dB,E&<=^LHV
J5;e8aA]K9EY:.R^K@c.-?[@dB3UEC-XNDS7.TQ9B8&2><a58S+X/E4?6]OLNg3)
aMQXeHfF9H4YM0fORb\6&\F#J6,;ODEOO#CG@,D8>e;P]T=PRK/f0LeLVY-CJ+G5
<Z1(#X#A;7d+(XA9QF+6#1RB@+=?M@B/QFFNGH-N0bf/g2LT16+5GR9BM=X\[Y-K
G7&N(f.((I9\R]YV?Fc=L1Y^;TdATY:[HX2L--,3@SS+.3M@2E:,?)_3_FfdP8U1
ZM1HTS]YLdbW=TUH?(/9NQZN_?>-K28WE(M9C+1/I&8-3/&^Kd=H(e(K-MU8JDA?
Y)c8abRd+/d.6N1S_.H,6N0KD2b>F+ScN^?@B4TG=F(AZH24QaQSaJb-C[\NWF&\
(3SM&PS70^X>1)=+P.O?R@[;)D7@Q].KGZU6?/CQI287/H3W5)EYf+V\QPXS)KZ_
WZ3CNc<cEL,Bd,)Z>f+[\M&3-R)]gO+2@cGI&aV3F=AF[1XP2Y8d6?UG567O_gAb
-DRSU;]a[bJO5T+6@4/R7YJ:Q+^[?afSI#SFAW_Q8U.c[-4SU@>Ye_#IdZK[e->_
=X_g#d15D,)XE&J6=:d86>\I(9HPW]F,,?MTBCXSc5=M)<VY_[7XODXScZcc[[@8
cGc8eK,W61g69gOP-^ZB&A=46BHc/4+Mec?)XA-Q0Y.0b@RSVf:/H:R[LG6gJa3Q
5cO[(K2eC)(U+D1CF8/dG#:CTG-AIQO0P5R=TV?\_BB@?@MNfc1B)>]?bZ=<dUU-
;/baOA&G+U<JT>?3>(cC4MQ<cN2=].NC##W:=:,>D)^Lb6\AM8NL[3=G;X@LK,Q1
Y0);QC6LMV[1;_>F,4P;AL1&SU9AIc]LVJ/5a)Vd4a>R=T))<:^&ME>aX,[bEG=C
7.F#MO[.37FUQY5bKWDde8Z(&F@;);g:QP<QPTXc3NXZVN^JX:LBG;T+=Q(fX1:Q
Z[?@J[.PWJ[3\,\#TVK]D/2TYR+O#4H:XFB(]fRfYX3,[+X.[N[8,O:9EB)+77_<
/b+THNJ;T9EVS]3&WgX0OI,=D[]?;FA[EG#IP]/R8_b>96?B1LU7ZM<S[G1;7f\c
fB5,DTWQB:cI&6GH.d:1Z#6XT#RBGKC44[dI(fbAP]3eBX6#Z>H]SQKeDQ=8Y[9D
9aBFOSQ]K^4Ve2MLNBXKdX#OcF<W//bXg,4Hbb58b+gXSZKH]ULU:.)VS-IFD\F?
53X>(4YOac\>S0]8KeISL^YBKd)BHa,E:ME/(Q90H[e?)F[K9A&5=816:)^VIK&3
)Pc5+=bQQJ^-71Ve86cL&(IKZ8A+,W9.C&BA)d5Hfg\Z(&54)[QN]TIU9W0Q^A80
HYXK9MZMZf4Q&_Z/D)#2L1].D(091]Tb7W=c[C0V#c<2^ON5:M+:]E/E(=Y)Pa_b
I1MB_UXQ[A:7TNg4fa[WZD7JO>XL=fPASYJC0=)9A_dG4RA3ABU.RfUWX(V#QE6]
=6Z3&H/&ISDL0D5VVT##a)R7f<FZ),;C2+[#Ge14eEK2-^?\O,a49/QdYS_B&2X-
V;6V;g0R&?eXO,M9+Pc6g>[]f[-VSZ=,^aW6V/-(NR?@VaY/=f[VT,bJ/\X,bOP/
/C@F6f9#3f[/(&;:BRI,W5.U#cK3NIJ&XB71LZeaTVY>7L32.P#,NBd_^a:<3KeE
,>HB0?7D>2N7Vg[,[LP_VO9#8:V3SFV4^;HdO8F1fU__YPSQ#@NIc9ZcF(7OcK6a
g1P_(W=C,JW3b7JY1aRHH>4[@M&\ZHL9/NLa6g3MJ(1;Y55G6-QeJGZOfD_HIX6>
NJZY8YYfUH8FGZ_@;&6+EI<]U<7MI?;L9>L5ZJ=,^Lb_aT8?[14_ObTH(UK6XEFL
4^3TL?<c+J#UYf,]Z..Z^P^XOHU^S2Lc:DK4RPMT(CO/34456H,.0N&.3)9#H(Na
(COHJ=:K9WXR?b.OKXPF@WW4:5RCXY<a+=59eYNcU2N9.A-;JF4Tc^>I[Ve&#,(d
M9NXY9QM&;=>F0\H<aRSPB6O7:fW&:9-&4gee45Ba>3@S=/?@AW(=)0d_HO[,\/G
d.,F&+0HWVMf&V#EC6MZ._c[d3[3aS30c7+J-?KKYR@)D1=N6<2.^[efGD#:GW99
@U6B/<.NSC.JQM@9.X&a:<3TFFWOL,MYU=4L8K\:OVQfF3O5CW]Ib#?.;2Xb#68b
A\<L_BF0>@RO-QR2N;N]WdC+cd;^9R>ed)Q_ZD\+PCd:g<d=P.AfRJ#INPZ[gN5S
DM9<4[M3a[D:bN,]DL7@@4X2(?6E#7=AN,6J@QN6<8Q^+<_/<.&0_D7e/NFX,;:T
aM\,OaKN;&,W:L94C&K9cbFF;HZ?,<4??2UO9&BY,)VRKQUJBGfgR=FCgN9^2L>>
C=3<01[]KZNX#:F(/L<0FQQF.34N>O6X2E)NJLC]]^eA@=;)K4dQ5DV,0W?RG#&M
7PY+_[Y.f;;M=Lg1dQAYA(BTIYSS3Vf.MNf07Yd:V#P6X3I/EggaC9a]0+gO=II\
K+CXTK7</=a:24I9cV&WRDWNZH/<8]F<K\LU@TNXHSfGAMXAH71;dY0/-\g^.@\/
[DAR0QU.S\YScf_9/+V^C\G<]??c109X07;#E3B3&UZ-Q1T74?U2]1<-\Y^(X07N
C_<V09D=e(?9?eE.J[U)WU[@Wg,9=,Gb;](2g)SZOT([K9,3F.O96(+=/PBXf&/=
eZF5F_8F=W9fYK)SWM:32I#LQG[>[;.PZ)=UVb4<E^>J(/\;J6T\/#5C[G1L#KU^
DKScSIYB7UbQ++@]L)X[#NYZ/]\@3.5M8[gJA@Za;Z>FH[)^MJ549CZ3^ffO)^KV
L2@)VWJA)d,&D2JUDZ=VMU^F=]=D&^/P838>>fGI@T9Id4(ZQ(#c<d^REc]W@b80
9c6G.]H9BVd3[A/E976([R;8@[dN6,7aO;URJ8=09\aA-5V9M:Z-R3b9L,?)aB2>
W3J=5N/38ODK^EfHT)GdG_XWN;?^KfdAA?M9PS4@Y3V?HP#Z>d93e((cL[99JF_\
#R3GL-V_DXGZYHL4Z-.UB4QgaY=W)]bd?ERS2A8YF@N_O-6^DMR[G_H]I+ff@J2B
A(bYb<]R)52&,DMIWB0YAbDGXZ1CXJ6BS+VZ@PAZ+O,@ZbPHJ._dTCB@6G]G:1d9
b@gX^2>+U1(LCgYKTJ(A<e8Z?c\Ta7eUOeG0=?-[HP@9;C@c?4Q=H#ZG3F4MV_L>
cAQ:c.1.QY9T1O65N[PF/,ONC(5<4dJGYPC/NC^eH(4BXE<V7I1#H&TM?1#:#6EY
JJ>]\T(0474>3F+?34UW8><:&-51c:DQ@R@e^dQ)X]96Fg\),#<3dA^34N(9/F.X
SCS9C/]E#D/41A(5ZdB\C73:@@=E1YC:F2QcEdG,fd3ESZKFG/(?NFU4Tdf?V+T)
+M/CI)\5B^EYJK=0/2[9IVB-6UQI3@R\F?C9WF5_Z-_S&#A;/+U:OYCeB+;+(=a\
XO[SFPO<#E&8=)1LIU82#Xb_3Z6]a9dTgSK]DN>L-1+CIGSc];F0CMa2J#3bADBH
KUGROZ4<ECTcTR;H#PW9MfG/Pg<De36S,L8UfVQ=cA;)g_.M]:BcR^-EME<+9cHD
4.X;AFH_Mb]?U)4fF3/,QU:[7())Y+S@g81?P]HAOZ7495SIgP9)(gNU;#^I0\E/
d:>\LKe3f9G=[HQgT&M;;U-]d#:?DC)eGc/9NKf/;&^;\82Y2^=?bAJDSgaJ0g1U
(OeK-0eD@<#K6JV/_aW[^.^MEf4>YIIJ_H.TD3a?69SYD:QZK9PSN2T+GBc?NW-S
S,3OJ<e@dCbHKZa=(6S.S28UeAbRRVQY;A\&WDRK0DXOMQ&Ee./d7WA4_B+/P@N<
JP&^4e?AI@1T<S#8b).=Gd]/ePSF_039Wg-_g8U2)\>5IF/B,K17c7DR-6dUKET+
I\JV1_>-&O?<ZUJ0eKbEB?7d9I:c\9HbWK652Pa:+/V#41.aU\PZ1(7+MCZ5MD\;
:8+?b&Tg+S+SRM@eR[(NYHX10--L-8S=(Q=N1KPeW)&KB^cS5c#]27R#7T=aEGd[
?6(Z9V\Z1GNJOT#9Gg>RRG5Rc@+,5NbY(e<T233E2d+)P0MVLb#[]9F@T>0;10W@
(G#17=I-9QP#>E8UOJKDE+Y(W3[&+?ZeOA_-fXYd_1=>+B)[-5/EP^W:6:IZ^=0B
R30TS)aaII?J2(N4e./L)\aNYLbX7cMEY=A<.d(O#M1:(OT#CUV4aP+f;]@<c5@]
[b7:43+G<F2-(:OG@F1K;E7Re.3Q;YWJP)>S4YTPL@XB2(63)AB+LO)1^GOg:W^O
g_GCbAPP\Y.Qa\1f].aCO?OUBeaU4@88,a<E]C[YaW.C_K@=\9b2SFQ+P?Z@V5:[
\FV+_N(;O[A3&eL2>T\&6SO.@JU6G#?;ESBR?VbA4d3V;&]3,bL69,NdbN+b]P)e
38BQdSX?G=c4Z1;4>?SMIS9LODa#?)A7W=E(IJ8]>E;/90?IMA6LC@FBJ#<4Yg[V
3]3RY3=Z^515E/D)J,;J=09,9-NUTR&aIWM[1Q)1]N>VVaa<_^UL3G4R.J2PI8)R
=?&@/BcTQKR0;.6E&LT=[(<_=CP1=9Y<IZFOVgN=?:Mc0PPcN2V_HA\TV]2M-H0N
>4OE@^OF)&3^[caAcf<bFUC9NHTE:@#gUZY,9OK-cba[@aAXWP-V+D>KX6^L^,_1
g0ES0W43IJ&/d;K+N(R[c1aW:J9WJc^K6;7J-?62T=c;\E9SI_Z6LNFK3,,.8[de
N3A.M:V?=Dg4U)5[@R#IGY1AfW\&[Oa3X3)OJXU(_#NE9#g55+/IU^Gg/DR,P-Qd
>OHb>4/#U.O([d7;BJ)f:4#gN\d:#c7F46eM2;^3]JDW&P.dcUaf.<\-HPH?BU>U
ZJ\c:@cFUICW7SY@0PR;Q4VO7.25]-VKNF.^\bWa-GC2,Qe1_.ZVg80a(g7EBYSD
TEHcW<B4,Q4Y+Z-.@_[:X=QJbF#;6C(CS/S@S@H<^OP;g0141g9dggI2#N+KE3@X
[6PQg<P&cf/HK^/;>-7dGMaS<YEcFdVa84T5Y&O.3g5D9C2QQ?,Y8IZ9GI+efK#_
)[A\/G-@NBB6H/f[8dUL/=952QALHOR5F#g8ST3A2RKLNf=T8,aO2,ORK6(&XIW6
<7a1)&Zg8edQgRafR^?YMI#_Q91STcX#ePdE=D^MK<=,e(-?6fCK>[OM-<+T#+\F
UAgdR]5&C;+HV?_)]&DeN/e_<E>>VJ1JU<?(>Ge?.QS6J1O4&PI:&)F>_N];)<9[
ENOgEPUUd]2C:GQECCaKbc4c0L/_dGcc1)GI69;UL6C&H<.KZ?PZ25MUV\@N#-GD
2G\7XQ_MV8B,I;-ZBK9NCcQCbf2<IL<485U9S_KD]M9P+VXD@3HI[0B_+B?=5EgQ
4MbOX\QeJbZ/N5Q4X&c(TN1TbfJIZ+1R>7N51&JGg\@bER3M<5<4DYJBRPK[Nd8Z
7JKPMAR,UTOa@22+Y7G^42.gC1OW:&&<Y:cA7#-7P]X#<K=f#_4+=NUOMF<U;d1H
V@+T2dX:d3B(]&R=ZGBTVY1=I(aT-/IH1G9ME@RfXaG_YXa>7SUP+KTM6G:>f#\R
g9#]9+fFZ^dK,V8XZ9M\1O+54bY++Qa56W>S,1-7OTD[BEaI-g(+X(L=Y8RQ+60-
Z//1Jc6CEb?SfF\2F9dE2O8FeFC.PI6YO]FF7RSMV;gJ_/PCb7N??Oeg/V]1<DWO
9R1K#O2d\(5J/\R51C31O[S[f_5&0Y;4MI^Z)&b9R]=Me&O]:f01/GNR-S@dYVgE
_XU^IWaY]Ca?A086+3^GK\TZH.;D&FAeP\B+.Q5[<@1d2[_d^6/BEHQAO,Z<74]V
NO-)WH/6AVY9H3)2H9X6Wg)IaDaCOc,<O#d&W+K)fF4@=[CHE.gRNVMGKWZe_CLR
EGE1KcI&\9F8L<b_-4JH\OdR=P,#O)g.>B0CWD4G,-UY55?O46c-#SXZ;^-EDT:@
TPc:TR:X0XFRYE=1]2ROF)FHeF<HQY_G],0JCZKX&#YE7()WIXLMSa.#]3/B(TNc
9H.<IN&W\/R/:D#F9(QV&fB62T0.baB1-DL^:,Y9d=GD[M793I4?OG=N<U3=VQ4A
[]Y,43aU)eN5G<HA@+,,58HT=[-LW;3/QY,AD+LD9^-WYY/#29TgWP3X#OIWX[]A
LR9eJ=E+C9gD<@<c.\f8PJe\(LM@9AV8NS7GQ&(>[7L.0@@cG65JaELT:^@=Q3f)
]1(\ZE:;b(#MDHaUB&cg\L^,8-(=;C.RL.?OD)5;6#]8:=#g.+Q^,A]S)C4+a6S#
(]e],=5Ue&^;fd^c<33g(HK[/&f2[K#69_\1Y__PMZDO/ZNQKH6/LMRQMg27VR/E
?e&(WW0I8fXQ-Y8F7N9Iaa:Y5LHEQ+XA6,<9QX#0/35V@1AF\a\C:?cN&1/K248C
]bOLX6T_0RO5#I0G8C06fI;YABQ0G=@4(cZ.^.HYI4;1(=c8d\H-dA.HP914VW<W
^&JEZ_AW#c0JGP^@Y,M8V@Z50LaONfFZH2egSbID\09BK1SD:7:_^@I]7ANM(;B4
+1bEc3LTdbOf7UCN2L/\Xe0bO>]<6^:,&XaX;:URW>D98T7U-8&8(FaCQVM7A<)G
9_>()=a1_#G81Td+K=C4N5LEB_&(Q>dUTYOWRRJA,)Ob@9\^c9cTOgUH;<,R9V.+
+Pc?-?:/>]aVJC;SZbHCV?H0>&WT(Y=SJBNAO.eG)0gE]#TbN+T\.M81LIX?P903
SK6Mf2eHN\#_+H^I9,F1]/5^&LF=-g8U+9PY\QJ._M(?+>(LX:V5>+V/=+PIYI@_
FT9106XJA9aVU?;cGb+EQg3S_/^@RMD;X)5D1#131XY<14I1IVAW#bFKRf8AT;eK
_[>_cTYM^4:(W^9b==aS);GV81fS_gLKL149:0/[]a>P,_<X&bDQFN53;fd,ef]#
BG9?aSMH+CX#)7bDSD-H2D?C#)D=RH(#/TDCAI5Kf]H,/c89]fbV<D_JDcSdR9bd
,6YM_^)/:4Q:;K\3LL/,6;8,Ke]b#-J(c\>A7]U@,?V;0Tb8&RR5)WCHT);T6?N2
NbIT?7S#S,,.c9[8LLb=20UC0/WPId)RL7<;7UVAa=77>94[<@.P=^7G&+0?d=>;
XY5)\JP([G5KH0:#bP(ON6N,#?Z[+g.WH+(<bBOf(HMZV:NI0NHC.(CXQ9X@Z&:b
W7K]g(>U&.5\H#KQAIdJ#5-=WK+6SFKYLU4f)\T(FI@]#1]8U4SDXc00RG286T1d
?:ZL@Q\\F=.38(IC>)RgF?J4CeA[?a]W)BT\PIMS;AS<ND^-PETKaT;\XYE6V^QO
2XDP3B(cH2QEgZ+ggdbJ-S5\:1b>M_NF8Q-/+CX-?IEO;&&PVb_5YVK5+a(8-IT#
YEL8UL?f+HQ<-YL)AZYbdDgdZG-O(]9A]9-M.deSLF>0]OYC#&IQR#ZdgVdI/b?W
c[CZ=aMcY6WP9/2b-:=QV8MK]+ZRdVd1+A#Ua4\C.P()cQ=^;9ASc5)K)bJ#4C3O
=TU/&B>90\MR8AB,4f,IeHG2C2Y?S<Fa2QcbbC\4c&Y?f<agDRP8;U?Q4;O>^&Pe
LM5aW]R3Z.)[X0.&\(a(=>5?WT)>9R\4Tg#P_9&NZ/_+EeS@@KgRNJI:\f9)E)9U
a;#9-daQ?&@+-M>168+G^\.fN_>f0W:be>:2J#AWA=E?([T9>:.S;TS?bGeQJU7#
C28P_(dZ])E=&?\\\[J#T/g=^Ne-7[X78>3d+QaMdZVCJAPG=Y6B+2d4GB.YCX+2
)Q3;d9.Z)_:=9S6M+),a<)&?.QHcG.?=I[/-\6KPBV8e51O2Yf2^QU_()W9/TINP
Me<XMFZ19:)B/Zc^O&.&FEU=7^V0.=cRIQ69CESI,=B9bR4]>?DfR9Cc2]V;93W=
9e1?S_YX5gWeZ+7,>ecV:RP.dPGRQ5JaW8NDAK(EQJ9&dC/^<eANFdg=VAY2\7Re
41VE6>;UE_R[=;^YY+]533OdGN-<WU:d^9L8I/=eAD50?<f6MPf-.f]V)G/cg+?A
X6:2?OIY@8],F@F^-Jc,\<<ge\F,L=#AYa5\9^b\]@??4b4f:Mb2#NXHe-,eX#6_
RRIF&a97NU>X0[#E?Y(Qa#:OXS]_Xda-<EN1]1/2PfPT5UT?SGA]6+D[9Ad15A+I
MMM#5f[\FaaD<[9?Q4bXS(\(b;[HXa=5;\AF=2/EVT,b767O2+dRIcMXA3R3/#M1
CeR^IMU&J&<[1gKVYC&W3@Ce(&R)]]/&;TO0/9cL,bWeSVc,De6Ca0Wa<aaVd25@
CcAafUM)VOSGP<CfM0S^JC[249@-F>BfXcT@##d:AJNH)W,CP@.,-9M7SgKFGE/<
()aggJ&LQeI,b?RK)F3fG=/J<9B&RQE97U>AY-^f/_F,0)CA49,a::BW1II)U#M8
.+@eI(E2?_\a&e)J^#J5f(af1&,,S\9\]0ABK@KD3IQ#V4K:a8P22U\6E,/AS?7;
+UP[02&1,RM]G\>7I=-@FE@MUELE\&^G1QTSMU3/TKL?OH;gAeE>^/M3Ic<ZHP#?
FXF]=.03R>bf_)MSWH[;8_gR&g42W:0C;RXf1c?3YJ3@O5J[1)0aFX<-T6-^c?;a
\11e]IAfS<WT1LD.S@>2+9Kf>FSGMHTK5HGFN9fR)+HYe3_EYTOQ9Cb5O.LRS;J;
eVW;,/(/.S/#gcXR@.a#U>[U2A2>Hc6B;OHI1^8a^?)Fe_8IPSLA61/Y7cE;gaKO
gffA)K&UQ=H\><(;M\>C;05cABdeB(Lg9.ZE&WMe]B(5+(R0@FC?^EeRW(S/_I\K
^5113bDPF.=F;&<U3RLfIF:RI]_&8OXU8E684L3JQaMJBT:G(DV58B[aE1.YS[ec
XN.<DDYXR)[RIeQd]6,:5M5YCBWQa/R4MJPGAE4+J_M7gHT3T[6g<8B+>e2U>aL9
dQZd>0R=eY8_B7b0TUYG=CZOd+P]8#)0B(:UeF4g)^2]Q?N8O,7cNTSO(V16XL;6
b5KFM(CW_<PGAZc[C]L>HOWC_(VBR^WXAM@LLMWg,JFY3IDgc6&(=I413fZ?9IO\
;_>0:?EFCIbO4NJ-K836EY2);c1GW(.7FJ8GBTQ8#a=[BP]/dSVXM@JX7N3]).TE
]PUG4>HW;<&Sc95Y3W/836>=AH(2S,_K:M8c&NWcL>7S4IB(C^)-/ZDAZALY6X2f
?Q^a(JJC1a+U=g&I18bC);B6]J6B;G684)Y<6YC+;[AI;@I#5,(-H98<IV>CE3^H
O0,WJUg0@+R(KLHgX)TVfHE>-<3a[/#S@9TK=Y4[D,BC(+=IJ/2?=d#/?;W+&PZZ
f7ba:XPe@2_7TO]Y6A8F.F=),47#17)T#5gMC2D_g1e-8F^T6E549=\KVJV7fO#X
T3BSIOea--OJ)9>1(+&?X9&>=aVcJEYS(=gI2NGZf[-)6&:,BNggc<GF<S&cKW/D
;E\Z[Cc51D4eBbY\7#>+4]bY-#4cBUO/)gAN56R)gIF[X-:Rb4),f\+\4b+ec:@5
[]9X^C<]H7R4fHDYJPZF_K?e4TQS08._YW/J;C.Ug_KY.=:)\-+X2Z4K+XUS[8H^
1dF1CM5I6B6g-.\CR&@K&V.cCL<2d+[PSGE_M;Sf,M=-&2VIcW^OM>_7f;@K&F9#
7ZSPH)E]eXL2eGND<1eO9K+<IOJC+ZaH>E_-N-4NZIf0IXPQXBg;9[T#CYD0R&Y4
#+V.RZ5,4f\8EMS2Z=4IEa9#:@[LT)HNI87->e^SU\[,PJDJ2Ic7,3YE1Q9-3_Z+
/BdAE3W01]SeQ=;(<f<HSZ&f/PXGe.ZMa0F?8d6<JB8FSIJ7WWbAZ?VUQF=g0JPM
f8g)c@3K?6ZLJ<9Fg6#Y.3&f?)QG/=_/K)cC+?0ZR5AB9)6ZX\@W\A7KQ:.1BQdA
W4^+U?)M]J4+H+MN#._]G9E1WEL=U0;7J]g(14+6d0Wc>=fCTd\gL)cGSVfFRXRA
#Y,RQdMf-U6MRMSF^:f[fAQ37O]fZ?7:_(71e#=LcD:IZ&8#>E4OLVbZ8MYbT?UZ
g#P4dfL#;=TdL8;7HM>:(?MD3gQe40[_AHG1Q3G74:-e?FeVEP4H,T#)JM\/9JP<
>84_HQ221>a4^L[=.[+G@KA<H,<(H77d@-Sb7I#6A\XDaGcR-e#g4ANc5M\+QL-.
e4J(]IO((<@U\[0@3?I<=Y]Wb?eI4FNd0N-eE#?^-1O(8Y=,-H?:@)H)9egXc\47
3M=O940Nf7&G@ON/=2bDH8?BZ]H=1=,S\]\,3>IV(8X#cFC[d^W/SROUW5HF;]B6
5#.297DAZ(#=,eQ)CISEfWPBcA8cD@bP;59]C^HN6M12V]eeSXCLV=OXHD7P19?C
P-A?;QHQD\D[-2deZdV14RQ3a@1@cR4b1FC/=TF0W)a_[P:HBM/DPbbcgXP3DbS\
V+(7-/0b_-)99/3]F)VMd=K>7DHa]DL1c@7K1d4W=f=OI]/]POW-QK7EgQgVA@R\
XX?G[N=9MZ[X#=,cf1O@H89)\dAQ3S0=&Xa#C0.&XY#H2FQB;-a;R3ZKT@K[>5:(
TX^\d#Xd32NY6JO,B-DI-Bg8fH^K:]8J1[V+9-&(CAe-efY+cLY&I913b#)>AJ./
O,_P,O.Sg)Y+-?,M0FX=,9)C.f@Zb#?>/6>2P+A[,U&O0R],^K@.Y]30=Wca-T8(
V,\5<@eFF7^G1Hf[I-QAMV:7.5=NP>JOOORX=;6K9MVM9YG\bZbb-]+I)05Jg?H1
W]26PP6Z-^HX(/I[/?N.d7-9\\-4X:4>>:K8X1]/0FU^]#eS>T1/79=@.c8H1;PD
;)KJG6U]R^:/=d@\HMd,8eG];7>X#)Ef0O)HHAA<K:VOPc]Z+<GRM,Z^/(M94X<A
#/9S:5d6?]>Ce3cLaK[6=;_]/AC(VN=GZ2WgG76J@WMSM^?<;:de1#)cOSJ\KUA6
&I@ENTWEfK2-?>K^,2a=f&&[[3G;&VU/UD2fE/g)#8f/0#b7Q\bg,Ud-0A]&T\)d
e[.P]P4gG[RA:g:I&2ZHN](1O8=2ME65,?&#A8PKdeGU,W4I(cFgaC5;P)/<^ZXb
8J;Z[9J3\;G.-]GF?Ic-]EOHOPAU6N48=Q=&=\8UAU&d7VUL8_A;F6H9Ge?63FVF
4QI>_gU\gB\:D6L#UX7BcW1ZMBD[?#TB<b>W-g>CEg@dd?AYca31[TfKQd/9(=+C
#?H0RUdaY8J.9ef=???e+RCcg(Ge>J^Ae#8/M<Eb3Id@@7_0EPQSTbEg0TIf;2/P
0fdMHT0Q.)P.D>N2e8WC6W<-O&S6/V:R\Zf7NATW@V-O/6)@#)KMOA3dV6]@.+5H
Z2N;H,aT>3Y+.C<;c.[N8UU1:]KdP7VTG4#,=D.Z\9gc([11-75-(3_K?0;6#,EM
&@1R+\KI(K(Z3L.M>)GX[0H4[@1#+;TTcP3(XKT0GAY.]8TQ]<+)8\EKN?<>O4P?
CHN67\-[YE&0?TB[/T2,GXF@K<cM.WS)^UD3NWG.)3JbIK?54.cg>d3Vf\0S.R@.
E6aUD2G>AHGC(]Y7Y/4FB\ZQNb+ITbf.M1E&VAA-Wc8SZN1R?;@)?#,##^.fP+=F
@:g+6GTUTHTPC4;NU\>;g<]UU<,QSRNE-G.V;J:feGT58IEeZ9+E_^b_Va7L3_9W
1H8ZS7L#3MKWe?&#Z\ga/^L5EPGKK7a<98MFa+0]ELK_4NDT;2KG,fE/Hc)9LGYf
7>XH&AZ3IV9E<_Z.;#9D8Q6C4PRQND7=0U9Nf>GAL(DVI&TRR8CRWL^@7Fc_^e)C
O=fR\eI:PA^:Cf#HT+X7&DY&0@-E836PP,R6__/1Wg7bP>9<&46c.X?5eG_d5KPC
:C)gePBM(P5SF4@#YDH99&R5DL&ZMYW9>C10^Hd_)#2Og,gNa5\6]4A&Q<V/]eA(
PEBe76K6Z_XK;aG8Ndc8X[S>b(++NB\^O>dW3)C]ZRK.#6+QY71/eV]KGd29\AXE
WW7?JY_BN@TcWdd9\/B3[>9+N/;@1(/a-SY(+@ZC.aU^bK7OWK2D<H5T/gW&1[.d
W#VK(]a,R-).+149A(33cg;54bWZ947KM@<BDQ0Q0#]7d/KWH?>1TQCY78R8:F2H
UG@&@Wd<:MS_8CX7cC2c7-(OZ#bM@ZF&5J3BSI?T0g6V>X2Ba]c4NSg>Ob9T9X=Q
5YGXOYK.5V;9eCa)6RQ57AgHZ(ECCeX9.O)#-J#R2;:,@&8;IHg1TNI[e-WS]4F:
BNKWaZ,#GB5WcO]3KUJ.HFaVS8X5cS)[1AL(H=K84X0eM7OFdQ.=KcLaD#J81B1Y
M[@;CO1\&43b&LTM@BE8b.J&[,-S[C^]ODD61TJH1.T=,;BR=YSgO[7VPV;7K+OK
a+?A?D8.3520^1UPbNF5c/Bd/;G.\DV)D,6>OX<\;7A8d1D)3;b22.#H&YJfK2&1
FG+W)6E;>CZ&eU,^f]6SB?6[KH8#>fR?2AY>3e7XL1V\B^W,#C]:_G7[.MT;94cb
J/@K&3.+KYdE_O.a,;@3>YcS;27R2gYA15VECM7BfYOT/M4(S83[,8[0,N\aCWC]
.:43S/JD3,Y^UDg\a[1\:R<F(G+&75W2c^)d@GR,W/YRH+T&_I]6#IdUC)VUJ][D
./1f6P-XCfWPRLY<D.IfE?4dWAS:MS^I9XUcSaK59WPBK_AOFfE^3P)F1K+Y&F?/
82LSfUGE01Z8)LJYYYTC@&:gSWFf@e\O/deVU?0Ob8&.g<2N[=I1XJebMX+QObYb
LCZE)G,g8<Q0+3aH;#.6O)I6E/J#TCeCSHcAdSQ@1_E;/_;.0]Q_QLgaXVQM\[18
B-=BE[f0O-@TBOQ&Q-152XK1+G6H>+FO5Q<&Bd^fA\Ma(3WK,8=58^U^^K,406g8
Z&JM(L0HeXdNgGII59dL_Of:c@.O>R<Z25;Wf<Q.6Y^5T^1gdX35AYX>U;LRY&JK
3>g-D^4)7.3MAXSG+,d/9R]C@?/39OJ4&=2VC&V4&_;WWD88H6IPUM(Add]6CCM:
>XU67DY3??7YD+Ad/A54:7Zb)EL9YdK20IG56.Ce&4#=XZLZFBG#&X>)^cD07/OH
Z_ET1c8_6b](,SKOaWb7=0Z]M&S7=@3d;:HNY^Q9,C8U;\_[23_#^93PI,,aRQQW
CH]YK]+_1EDT?B9EJD9bT?2A>edHeRY&;KA:/_O/;68Wd473CJ(R=Ab#X\+)-5X2
eWBb#=<;\H)CbU9K;D\[-_=/Wd/UYFSEWU\0&9)VcRZ11SN]O#@P,eCeT2I9WZ#N
6R1[c4MSG2Pf.T+[O##eM9C4gYXZXDWSC8b=?&NVJ6M2)e([Yg3f7Yb0VIF(ad8a
RaeCNg6D)I1_C[.I[0TL+0X)U//S/]&=F+/LX/YV<EY+8b&2a,<8>F,37d<_g6A<
bV=S>Z2NScF]E223X.9f]9K5A0&VJ-JDHDQ5E)eXcV,GTUB_(\&]PN6/UP7(^<0P
VQUJLBG+N9L?#[a38a/1?b424@8aRH9=Y>^C4VC.-,FH3[a<[U1(2]:@952VLbbV
c7@DfD3R(Z-9e<.de[=M[PL2aYE)>W)1M_G?a9J5@@_a-a1N4fVO573<Q;-6dC/#
62J[T/P_28b4eXI4K8&.13(D2(2U/W=a>;fBVIEZQZFA,;gdba0H\9TU2AXE,2,<
D0RC:6Id9b/9RWB:6]:5f]a_V_X<D6=NC-?X@e]@>3WT>3YHB)-94)#UKO;KD-/0
YB)W>G;V,A<3.BAQ2[])V7IY]B(U>:YfIZED2[0+@GG&J+g#_;LW\dNMIRCSU>b[
bQGAG?^O5@/FS@6D4QPG/AFM4_6bO75BTGf;_\#_30>P4g1()#X9JTIbeT>CCU\/
MEQ6e0[BQcDDCH;3OY<9g;?91GP-(a.^F>SX@@O3A]3V^H8,(H_#M/?A;##@>K_<
(#>ZVZ)TPCdd8fYJV_)\LTOZ0TMLP5W(>#agS_+0RKf0eFW=gV.d]:P7>CGDPf@c
+,bR;8-LeZ9b?dGU3W_AZAXMCH--MSdU-70-TY_&2;@BD+WW:CTR2SJGe-<9A;V^
X]O,N:MG00N<eHJ0DRD><R-&(H5;.&BIFDB]#)L0A<#D<^S63,Q_Q/8/d/XVR.:a
^JP=3EWf?HI(BGf4?D,FBO,R4SF/d?aO26bf]YP=MNGMCT(>0JY.4(A:\?MF(T/R
MM9_9?#?7D3+FM+CQE<:@B/bE5A.ef2T7+V\2gV6bV;M(LPYG1_<6dBFaCHef4N:
?RV.T2WO-<U&)_I@T;9G>YUMX7WfBTK>bUgbLY:Xf\G;/;E\cG:W#4-K0H2?^5^T
P4(6@54aN#b;:(,Mg;?Z)fFV+BFVV#-.B.aME37\\&Y#dDM5I;XW.G-dU8gK1QW3
T?eW;@8W,cDUC4MQ)@Rgg&]W6Vbf\W3MK.dWEDB;L(QURL6EE)_X+C]d+3XGCXBI
OD3Og)8TO13Ie-T[-a]6(T<?0MYA6;fC8/44^UaBC;SJZ]+>L#(f0VRZR8dR4.J1
DgdQJRC0\H(g@0-TaJ3G^XQ.LESIDIgVJTRE,=)3UO]MGP\W[b4)IOW6?YEI5+c)
0HQb\J0>4Z)\gO_:/YY5BZI8<L)G1E)f_&dacG6DG,PB2dg85M;SEgAF(,))CL^+
#f&e40M&A?,,)>AVPHPW3Vb4@];QA5H>8BJ=&#H:\63ANZ02-921(>,/S9LT#af&
Qg5C[C<MEDCf#^/S@+#KUH2V33/_g2bWK_d,)O0<SI.9/cCZS8a2M2B8+D41]0bg
/gY2(8KF]8:f_21YB;.Z9_2f+TK&012PB:3(P5V+N8XDTKPG7KeD_,O\+SQe6Sa-
HG\V)S/:<c.gQJYGS6+280WEV1ZObUM7\KCfRN\;2AM+e].6+Sa@Y<QYN0S5H=>(
Sf]MTUTR1OB<>;P=dgO--5a&):4C->-O_T]9Z<Z2SK\K/]9^<G2J_+&8<aS>Oe#-
c)->LYW:I#E2\g#KfOUfD>-(Z<^ee(9,Z/(PHLRLZ5W736,MHV([BB<3:\,59&]L
EI.@&S\fAAKF?/Qg1[&A/-M+2_W-b5@Nc/LN\F#_7=>_-1#Cf7Y_VM/)N;df9?HJ
SCVELYLP[12LMI>U:Lb/SceNW8IYa\CL(PMDFc.eX3#b^Q0VL74>0D]dO?B-aR_,
>65]P&5=B#:(eY]Uf0dM].-X.aYCHS0D>]/e5FS>PX-;)@V]XUfW0OB[&W0[JL8.
bPBI;4B;NIEgBdVQW?>BcaBE6GI@6+)+a>F[b@51SE7ET?JEBbFUFE&FeS8HdGJ)
E2J7e(]HIA;g,@/C<3b2427L,A3QD1?@b5,IL]&RT-4cNNd\,Lg1ef3/M++D,,A>
YcQTXg2ZDPDMAdY&Z0GYNJ>\TK3R#Yc5Wf+/WL:(3,[2)bGO=[^eJDRV7<3W@/IZ
PP.BOe=V#?M06UJ?A+),76VW1H-&H22#PE(X1e.[^AX<f-9Ff3<OE-J-@dKMAcCT
9A)BQI-Y@<5deZbX[FI,G6bE7&S4#]d[S@WZDMENDK-,&(L<&ac4FB1ZE(a[>J=P
]K_6D()L7V6/^.B/@?^=cc0WM-+\=E0S]0V-eWR<UIc?_(M3a_d_4a(U_@UH&LY7
YI-X-U@BL:g4,A,XXCL(O7O<P=S#Fa;;H0gWaG9P:;cJT1g[B@E#dX0.1,eV-ED(
\Wc(TZ7Wb9+ADAD]@<VRM\KJ6BEO9+F98XA;H5=@T#-6=UMK:R_Ig]Q[LYEKVTfF
S,:&P.[F^2ff>P(e[gO?WC?G4:EK1+gD?#Xf_c^K+dV^)J79Z\Z3I(Wg;PQgGOW<
2)GDGJRef_gI+BEP^^-[bD;\PL(S4IXKKcXP]#AI=I4F9(U3g;DIfNSc?S]6FSG,
.&TP(D/U62>+^>PaM67Tg/5XYf\D-^[+c^P=X#:Sf8?\Hb2Xc(H.;N\]fDUN6DHI
1F,M#07&&0Bg.MGUP@;(A6,;7CYe6]]DI[>WD2?cPaO:D+#Nff:#Ggb46OM4TW(Q
b/\:?MRf0E2[-IHSJ98&83L0c[f[+RM>YF6GM;bM[a>4\H&UA)DdSCD;d,0?)=f^
5B78K)94I@?FO-+</6@Bg4U\5:ZO1FM8:N0B3e1Kd^ef>feYTa(8XZG0VN5:EOR-
6T98KeEU3S_f.Q]@6&/d(8C?I@6]8D=+7B=(g-=188\(50gc^=SQZgYT9?R(f<Bd
TY:KFJKaDf0+1c-L]fBN8fYZc3>:M<AM/R)9VZ)M>&^L?UK5_5QX-EgRX;FJJZ@,
=4/d<3VeO<a9V/cY;MM,1MDQeE<=fT9]@,d(bY;Pb+A@618LK-Sc(:YK:D?6.cBg
WgSBQcbO:Xaf#6DCPA1\E-##0B?ee=P\gC]O=&dAF>,2PTZY7bL(1K-MR9:Aa0T)
_AZ4^aIaN&B0LR?8eKXVYK7]g;Z=?7OgE:6aAM&6/gZ0QL&dafd=3Jb4?G1)@)=I
F.H9&J2OQ2+<c;6X9U-bBY;X+>(@BCUF?]DbFA@G[JD8=,Wa0J.VXF@<SeA\1D_c
K\<2_IVZ1QX68DNW7PJ25DPPeW5AU78RV(?<54O57SOQBF)aM1X7(^b\P)#J9[L7
VC_Y]64EQ>C4ac<[+JJ#IX5A8ZGaSG<7A95+4P624+5XP5/aUA;AG(V06C2CFUTO
QFAEDE,=N)f:,Y:CP06M,]CGQ<Ag:-fVFY1dd?;:9G;^I[V+;AEN?6H:0a6@GWcJ
._;:\B:4UKcDV?Sf5<[8)@Oa&4-<:eYaW<+F]-#_XJdU=8(-2e)[Sa\JQ=.<_>X[
HF:6R9O-<MS\R8M9[5MMPO4ZT/GfK<+4gA2a&:5GS@T-[X@=55/Xe:7#3,P?&g^(
4#5]&BWO[8T9#[2BH,@Z\(,\:S2I:LT1K90-JGcBLE-R<7UFH4W#dcaQ;9TK<DAQ
c?L@0/_US-[H1\O\;eeDS;QG8HX4ZD&3cc(0f<A]S4&a)9DKe4N>R/V]1NgTQY1/
T@WbG9&?d96J?.R-JY?aYF907XaWPI-=-&d]MA4?bY^50Kb6N54dNZNO465JU/>;
Z6E7FLC7cbTY4-:[@3NR?49UUKGCTKc<:4JB,e5dXA[9O^/bY&HD>GBFGB9WYTF@
Q9WWaIbNPJ@_baR11G^VP2Nc<c+V_;O_)1.3IGD0?Cg=<F2&Md2W3a\--0I+c[^.
1M1CdC^,HPFc\UaMU<&YX@A+JPQ41T<NTaN#AbS^_,M5OUd=CfWc[c\(dfG2T^eU
Y>,aQP\XQaEIVG9_I-3#HVVWE)[PT>KR9+@ePGBOAI<W55Ag).:9VSSN5aA(N-<C
9ED.g-[HZ[TKNS-D[42#ZFI1A&b47b(,5H2V_ADKRRJ)=5^47gEXQP=/)WF560I7
3=f]()1AN1HWM/7F#GaB<@]ZT[]Pb##J1@;YL2d9Cf]\a&:M[f&=cef)1C>Eb=bR
?M\bMNM;NfWcNIU[[C&)(G;>H_da&2_EVS@g[<LF5TJJe7Tgg6R]cO7@;cg4>TDB
Va>C3df\]eYSI9<;?;EXKWQdUC1>ID9T-3H<d=25,0-;)PE)C#:AQJO6cBeDGbTB
O7.HC\7#88R5.\C/RB]f7U+^&)c?/G9cEa49Q:IHL4QPXL1=d>M#M8geKYccTJO#
D=.P88MRa=9/C=(W]cd5>JJf.:IWP9AE)CC+.ENOKV2[V,C>aF29bD+a-JM),2#R
G,Y9AXR@8:/a4b1DJ8dE:,+cP:0H>_GJQaBAgA,NZc(D;>bA5V-7Wg&f>/J]RW9/
c+Fda9E<=FRE9-6O?5(b<MZ=_+4TVD8B>gI5=YO5&;J(W+4(+d@1U:c9UW(X9L1&
Lb)AK69c?e[UJK-,HHP)V2^BJ+XTJB)T7USFJ#,bWcS9>9M&0.:U_3H=f\#AFIUX
WU9FS(9gfeC?T/.OHHJP2;J@W7,:SN+9/JHMHVX2+[gR\4)XYA6HWC0aX0Q#K+I,
^<0\AFP1ZgJL6BgV7]cWXRK^;NVF;cf/;0\S89S7-&5D=8LHN7ZFU-K+/#:?]Y0D
,bUEQH4./@:-CEcRCDc5:^HW6YR17Vc5F)PQd:e,WW8:0=I\1K>;<#7O32<J7KBQ
dZF+>^CE?]T-=@YYM24YJ9ZMd;FM:BYfW\+.gFCC@)R>XeRBTVRN3W?H,MLU;E=.
[F2:0ROQ9YPb<=KQRF4VcfUD;PSQf/91Y:-/=+X-0&+@WNQPJL/[?aa3F]EXV5&c
NNMd]e4;P2f#fbG2F:^a;Hgd6Ld._):.M[#JM,f5489-2]d)S>CH6JCOJAO)61S7
c+7WE&e]e];<]F8bM8R+9@_TZY)ag9,19b/D-@,RYT;/6WDGH4Fg2gMe,0RU;WR5
0;U>)+gLT]:T78F0bF4Re:&)FcU-TaeeEZ(+_X[<+BbO9Xd>LN#,T?>F(8fQ(]2+
f(2C(_LX#EcCAAAeM)19A33#QU+ZOc7F]KcB\1b&5NE]DcP&b6FXF3V=(QGO.M2=
P[2N/<REDL]FK?NR;&e&X=&[,-H_D(BKZ2FfJ54DQM_37H[7M9\dY[\9ENA@D/Rc
c?fTPf)@SGN4Fc5Z0b>Af,=Z<4&XI?+[V6:Y=eg.d&f+T.Lf.>9cgM,#[TJ<(&aO
JNLMSY,+8eB_2UD6[(^.5)#X9]N[N:)<gWRfcP38B=CcD7YBIOQ05Xe/9HNOM:Oc
<UYYMMZfJW\J4N^SQU+Ia@OeH3#1Qa<K<XCQCb8#,P4,TOXM\1+SAW5<HEUW^CJ2
K7N#T8aIV++SW2PVVa],J25Z?f^:ZSb7L03R-[VP,@)GQ(CREP(8/a]NJ/a/75He
?MQH/E1>RcA;&.FAVc(2RR-<P>V4K1CR#d6e6<bBMW-.<MU/6VF5[.HW,;Tf+BRd
_1W_[8/:S.@_G>];-8PCTZ7Kc^4UOLA2];#gKggHSe]<(\/SGGJWQT38OeGb^f(P
2I^6Kc7H/MA<00J8\>Ed>eE/cQ-?(\2B>/M3)/,OI?FP18F0->WIbO?g]<fQC4P4
^N.T&3IEE-]U\CRc0geaZ=/ODX@-I,QbP7b\]YD=N6>@:DL58EI)F3a8Gb9df?TB
[<,BC7JBXJ68+D=]=EJ7^C1f8<SG0+.eH5H=RS=E@A/53N22(]3?4\dYeaHRF3Z#
L-3K(0B#85ORa#1G3<dg#I1HJeB(24#X5RI+Y-MHI,W:O]5S#C\Yd9D0MgGR13O1
>G<?P?HVBIVM4&UeX/63J&.a0#g,.S>:KKSYDG<REIXf2]aMR;1JI,FXU95/R2@Y
ZN71a:R76Q;X]@b56L;L2#^06]cG:6(,3;DO=+QNI9?(FQC6?:1AIN>=6DV.VgU^
+9dFPW)/R+Q9(\C3Xc+WI-&(cXaMfVI0EZ:TSdL-dROJZE@d?A_=8ACQYU;cgO=B
Zf2JS[V=P@JCNXb+@.bJ/;9ZV51^2C-R])?V)QGB2Pf\.Y9KVQ&ZJ,31][X#MH/G
0HHAIHPYBD_I1IeKV52?PE7B?GWT:AP+#7R<>-GLcTJAKU;+Cg_ME.ZfF4_B>2FA
T4TAW8b_EK:X1Q4.e&:QKE9A=,]6OSYVWH:\I?+5\,8NC4&d&Ya=63<Zc[Q\/3MM
Z4G.9AK96KW\8aD:&?:+bX@&YL1M+=O,eMR/aPQ<E_eMMNG\M<@aI/9g2>(gDfGF
QJJ)>\#1@,LQHKB+YFaXFf:FW9S.KcNXD;/5d+,DG]N();U]KJROWC_-WU_RW[10
&O7FEd_Jd>GVfKUe+Ua546.H4Z9dObb3EJ^M<?>P1YB(<>cR>N,3DN;&/ZP<.ZUZ
bTJ#8FE_eDZX2127WcM54;;Uf@=R/D,W[f3\(g<+B/VaEV2;003-UT#US/<)>/)1
Y^F>K:;FBd2>3J<O1G=cE=7B>12Je,N\BHP?I3V5W#6[B@[^FV,JIfM1=d?B,UZd
>9&b93B3PALRJ_eF[8VVZ4D?L&Wa>7[I_VPZKa;BN/&CTF]Da<_Z6\?K.c4Z<RCg
R6MQU8,)4Ud#W<7-HO)I99eQCd&Zg9N6TS6)_X1,+6aN9VTM7BLcW0(QgO-FU9\-
=B?\Gc15MNg:Xb=c[K7fCAHEU(LAA>OKLP#T@]4@A1\;3g3JCLT/7+f#bbDHbRBd
7T^S#&;YW>:bBdf@R[/J,3FV0QQ<<F<aaE^1I/If5Had<#S/(I#[05+Xe:7CM>S3
^DV3A[N3bQT(_AQEBB,^ME.g/-.K\XYP+9;3f?[U&9U,1FcUP3&+MeAd#O.W3J9,
U<9O+d[S0]f>(ed>#VO=;MHf;YLBd69YUKG2d.GTL33a;7HC>7ZK9Se&KL\-7X-8
ZFQZbQ4RBPQTHA#MI726.E\,b,?&MIc#A>.9BDD)bS8HfLX]GeSQe&>I>IKD6<1\
-W=J)=VLWUb@]7#-d2M[PB)Ob^V^:E-@#,67O@T0G955@Q4;CM:N[NL#20^g=(3;
_b9>TDS?=OceMY/TdNX.84LC\&I+&1([f_?5C-4MR?YBbCN/:Gc_FM?\3<IYP?F+
ZN/B.DTGI,.=PJ+3U0,[B7b?]C28KAe22JQ.L6D&\@]gQ/]2KbUTD>\>Xa&2g:HF
M19TA1-gKU31B&=6>OYf1;(1e[W6V2OY_\BaO;5gWRe0>Y9\(D+bP&edD=@@#H,(
77N>53TQ-L)0@FX6PbQC_WSRKY;.>P^=PH8?>[)T)NVK-?c@@^3OWT@T&V7gU:1f
dZ.#(VA@g+3d)-A97D)?.HF&LffZB]C+FeGT3J=4G1M6Cf;R?IX7TbBI5V6W@YFI
=91^e7U15G4:L>3cbP/W)_4GQ<A<>CQ1LLTGAcHR&,HcXI(e8f)&8FeDW9CVd_UV
A(Wc5,._>e,GP(,;&29A->/#N_]Y,@:J9<#C<JR,K?_-?SA[^Q[?(9_?I\9-5O1:
>/M2OYQND=TV.97LfbJRH#_<>7IB;ZTN0P(2@E(&Z0<PN+G>YcIe]M7BPg;3;E.&
-VKGcA&3(5JdXB/,#I,=9NRBNH9AZ4KM+dRV2]5;&YW,U,3;VWG,dEF:NgC./M1J
#HMReY#]A5]LXNH^8&>AaDDeD?afGQST<S65=AS#H>OVFB2]EDYD.ZE,NY4EDf6I
G]_VVQDK<L[)\&e1T_Rb/WcKJ-,PccMIg+?1375#6BD^-DNQ>]QdVIO6JSg&W6bC
)FV@6PfK8G7b;<2R4aKM5H8,f[)<Y[E1@4\Z\]NJPTV.K7GaR/DRf3(UJ:@BSeQN
-+;Pd<dd,c:W.\J-L>C;+,3-aV3+9PNT&\7F<13&3_6gA.S@FJ+Y24)=BcCJ]<?S
(.D#+HceO;C(aB774,)DX(Zg_#::;-=6^(&UcJ>9.DJ58Aa)&?RN.>WTgb2V\EG+
O_]ORB#SV;4]+d4]R(D9=B_XO-0/T85H5RJ_VI-BF&+ZVTa9:6Ld_PCAC0[aHC[e
0DWfI(K&?Q8H,Oef(<RO[W.U/f4b1G;<<5aaeYCg+b\6@Y/c4/d&/;US1&R)1GS\
[<,3Z@GITCgW3FQ773653)SMBg5A4?afU>P+^D7?B(=B>Og5Q,<46882:52(L.=O
>AW?-H[?]Ae:d[GF#)3IZBA9B3=/<bB),Se/D,dM9WJEbIYJ(Z/=eb]?ZP#DY@NI
?Va#-H@LO6[P<C)gR=DI=B,X99OZ3X9TW8E?3(MTC?FeSNV99Q,Ef^VIf(O:,B)2
AG+&8]PJWTe-6&KUVO+f(aWObJB+[a;8S?Q?F<0MN=VA_Ic5EKO4O[.[?R2V#EXV
;d_BFMS0g8_Daf::S=-0;W\\1_I@CK/:Q6gI:+,^@RSJW0:4[g(IUf+7VFa1S4e/
ca3Q.FfUNcM7ERL#(?&:#7@dP(d:?(0>JdA06S48<Qe8?2&G7G^DO<26e_H;??2E
3_DAc4fJ]@D/,D5^<N4+A-OMP^gD]0cWf]SIKTVKeD?dH__L)DIdJ0=6,dRLM2Gd
5TcIJ(G,efA)C(8@bc1#_^#G,.&JHdJ8fG58FJ/HN>>&TZXNX@GF]3CMe;#A&,46
IE2aKd?US1XV3YV,KWBQ]D&gL8>LG=FQD5-XJ:35Z>I.#-?DLU(Q@-PQXE7U0_6[
0>T3+VgOQ#G@KVGX^_DVNTO+aZBQ9T97NcML1=9>GRE11M3cVC\JR_2-Q9f/6=3-
?Qae@R2D_DYWHHf<YUUX>()4.I;P:<?:(^Y-(BU^<YMC-[A[DbPH.NB[T=;@YC:^
Z<=H1RV/feKHM3572<2b(31<a1XJKBBa,^-NJ8NQ;Q4d(BAX-Y-2WQ@^V6Bf>682
@c.OVZ^^(:6YcY69XA,E5<M<J(GWW?@(4Q?5HBaX+W]C(3=aaegCR54@4MJPQ>A#
8LDR(9e^Q;N#B/5aNUa6D+13GDSH=+,8/2L:A2_T(UX/;X:^WFC\:,QM@;>GI=DI
ZLN?\4[>1FNFB\M9bKUKF=SF]))Jg-bd+=eVZXg2QFI1P4<X@Y#<4<GV=HX<A(XV
03Mcg<<#Af805.&-.J82C#cU79U1]P@IR1N5>a0BUgUI/+4JW(ZV(86#b:OX#IcK
\M1X:>ATOR_+>g7Y?JS,UX[;b&g2:.B=4_8&bBW,D)5;1:L)@0Q<PZW/D-,#V-(c
bcA@]SXZ4\RX8_FVMI01Wa6<^_G55(fWM?Qd>&d7>[LF^NS/Pb6&/.,0/Q#_7\9F
C)CR_0DfcMLFXb+bGN@WO#0b=b4#YV^NE6<6F<cMF7?=IfMP[Og\cF-HO-Wb[JF0
ZbQGf@V?2d;D6Y1M&_B;BX1THa3O.G?#0\C9K#(?JHIA:W4573P<aZ8-<Ifaad]Y
UB.G#^\@-LO,\Ud/7YO/QAJ:AIELV=M>/:<KFb3MY6EODSCT\H5:QV]dgNf+de]_
dM2D2c<K:IZB2T,,(5_Ge6NG-;[>MN+cd87L/CB3>H[;\NK,T?](g9W^(B.@00\T
1()[<bfLaWfA16O/:Y9R#,N:]WISK6&[W8bf&\X,HOPcS>:98GQP-O/=<dVS],K&
b[=QID0[0FHQ0\>=8:/;BXNZ2_^QeZLC)SAV_;PN45IB2g@/-:NJ4-:D?5Nc(N>D
FTe3aWZJ8TQ..RC[C6;K.O0.CUSD.JGU9?)5H-.U=\f>U>cPB\eDE?.G,=TVRcZ2
Q?+5<UAF:?gODEgHRNgA#3/=[D/GBKKGE>)abSgRcB^&a?g[-5PQW@34[#;Q(d-e
+,3/V\6]A,dHA5?7VgVPf@+#.M(ST@eM7[]Q9=U1<7K-TSC[^G)YA5Y_#3_4/P+L
(0PddR1V9CJ<;fYGYAeb@CKH0G>g85fd=FV0XcM-@O()MLF0:PX+E0X^BPXZgDX.
N]F9aNT+E,077X#DV-^S-RD?BO_U48RG\8@WQ_Q^K-I;/2U\3BW8f13W2b<QBY^>
Q-K@=T[M_+_UC#:]GG=6/EA-IU-#J<OES_[Mf#Q^0WB)0a.@)(P:1,G8BV)\PL_8
Z-,VTaa#TSPVSJRX8NdS5MI57]DcMcO#-UebJ-&fC@+a]+TAcG)>Ig.D>SU_\P:d
7S6;eSH(E(2B=20=D?MWc2g__C2S?9dgOKC#9(1@ZEU7,T]?;6OYg8:H7(]\86+P
e78f_<2I:b,,.]#KVUcBA4AQg#2+c<9&0[+I#?,#]d2ZQ@N?aY4b^b+.QS@4e.^9
E#2B/\YFSTFaC2>8Q2CBWUfDI146g(#cVYZ]Z(e_7GO;bcfNA+f;=TcW.#(SXM+,
Fa)RQ-SFT7+8<+U0\CO=Z3,7NCT8:9N;WW1K\MQE1:EDcW+aU2_IQOAB442;^IB2
]6fH^QG_FVXVJ43RUIfAW<Q6]F)Q1gVFe#U(aVO0_L&g5WTEQ:/1?M&>W67ARMaC
DH#16:]=@6MVG]YW(UUH2&S\_K:O#V;Q635(-OU6EbDdZO]O#S#4g<U?1<@HAHM#
.47)QM/+IR)P6a1<E^?U8H\VZL19I<SC77YFDVT72E2]-/c^RgGI:6bF+g4#9D_.
H95NDCH&(;LbI652,A=.6JKS9UgKP5Z^?GP]5.;d[R=I).38VfA]Q5E85(c31ZS/
)0[]D/^9MZJ91/=Sg^1/Y]bI8YdQI52gRVS[7&)c3D-Rg4D.<W_[@_J,?a\[WL#=
MA2QK4J1EI,76d>8#[C8)@9:P44P>6LJD^AZ838VP)5/N2/OED03aUY6:IZ,32II
bSP)LQGagga_B(gfJM-@09ZGR80OS(4BH8=U?+4==D90,d.:C>\Z#=C:9^MQ:#ZB
R:g_eW25=6_e2;Qc5\H-?B^#@+5&f79;^#_:VY@T9NGf]700<0)^S[.1(>;RD]A,
W3GZXV0J9JNP+MTE+R7DdMEKZS1PFDEA6GMM(9FWR8M9b^XaW_03fG7M9a953P;d
9F0RHHV541P#U2N,#d/5Jf(W\dA)L(a4_)JH.)<D]+=V4LEH_+XgQEA<F1^TVB/^
9Mf]#R4Z?=,&8I_6)6Tb@TF)4YE:W#^>1UZOF9GY4WMQG((D+)1;b(;Z^D6bO//?
FZDLEV=WI?aAF.-6A;A69R8Oe___<:=S9=[76JK;0dJG^3\384e)2FP6XFY]CKF[
5Ida3M._+J#Tg:9J\LW^+67ZBETfeP#eG387=R]d1c;L7fCN^#HX:K=WcMJT2VR5
c>7N\XXa^7S_7F]Z&P\7G;7O^W1+7\J-[cA]H]X,&@Jef0Y7#9A\IYR6AOKJ_&WZ
A>-B7JV.dE\X((4/U4/\MOc)J?)]RQY]=5RHK#DBQ5&([FG;@baGKR]2\6D<1^WE
__X^W15ZE>X#-]=Y^XZY1GeRSg9e_Y0FNgZdU1.eCL@8C#EdNG0EcTd@JPEE-:U1
^8@\=DXR>=&V,O.O,9OV,Cc^A0)N;Q?KS+36W3EebD?O]BR&IR7R6OU@EV:DC0B4
E?[=c+O7#-ZJ(>S(5_:1>D>8L:;/.UDE]M<B?NB71\4>/Kc#)D5R-<-TW?9^4/Lb
H<Wf?@IbXQGH1RU=7;:<+]3Lc2@X[:X2KObb[d-_S\WU8PAec8A0CGO-,(GC8T?(
c5J-4RF07LB;OF;>Hf=1AA>PJ)V[(3C?J2.M@PfbD2\?aOLe+I#V78aKaI+99D5I
2DE@8.]T-CY4aVBT;g5E10ScT_B&0dCEaaB:<g<ETcSdOIJSD1Vb<15>G@\75R].
3Zc9KJ&KROb7&7G]R,Og:3+)Tf<Z@MB;0+<P3VS#0+;Xef8(8U9/1@(?<IXR.<CS
J8e]+7Y#_<Kc16IF;#;+Cg1L#.OB^,3)(+)70U]@XB\c;<D3V?H>ID1-GV5,#KP/
]9?8FI1OW2K,gbJUD4A[>S.R/D4OMBHZY[G)]7)JAc51&76gDD[.JgU2:Hd)OJ)B
(&a\1WUa(:/=F=>?#cL]B[_20,Gg#[J3CPK]3#IA4gNd5&H44;Rd/&:f>1eUIU5D
8)8:OZ9^,)7<Y?E)@7SH?)6Z.MS8[7]a&dG+6&4^UBNefO\dHCF6Q.6e4I\8d,2Z
7-cRCg)8CQT=XDaR_]2#bb6LF_gK@G2V)Mf@#&F#[^2If.b&G)?50QdfQ05)?D]R
DGfZY#WQe1F+8\#^8#WW)cA=4dCZ-.U7;^gc\B4(K)>M=_).;S):7A9Y(Y2G[7(9
+G0SBZ2gPedA_?;<[bE_dLd<6MQ(?&Y3/6]7;&U3X7cC10TA0BG]E[+d(::-/&C[
g4IcH3U(+Id12D55=0EEUf;.a]RR+.0N<NPTNYDO-9c:VSS6+1De?QWJJ(?;9G;:
<)<fPL#EFB8(>?6L(.[f6)P)8U:5KFZI^H#K:VVTY\)PALD89VYN-9e=MOYfY,OU
Gg@&W#[.)ET&)0g&c<??N:FNBCU4K&H^-B8:(UX?CD6Pa?=L[B;V39?RKMIF0gQH
E1P5WC\=Z7+&E[LB_Z<L[73?LR9EW98OAdS>O,\9OA,MP^6?dLWf&J_gdd0O]aO^
+LC#?-4dJP]M<5:e[c_;)Q(.#Db><5X>36TZ@F9ZZ,=Kf]3cR>Q^bPRf_NH2[W>J
\4V@8<Ia&Ae1#\[)1KYOT-a/7GT_D6ZX-+@GbSLD@@[aZ/F:^2D#(;ZCL_7YbbUY
1W\@[@+-gFec)@QT/QL=NHD;DKDgQbA,bN@LW2[4&2cL[8R[S^J:aBc_US>X35#_
B?^\[5G[g]&c8@W9Z5)7ZE2Df=;IA_Z:,-R>;9&]\P4,=.OABgQW5RN?A9=,I)\F
IX2P^&#]/2.9&T4DAC;UZPI.8],ND:#Nf^C(a/2Z>,<,6NVQD9Zf1a=<QEa[FL[^
_ZOL62L/ZYRY9WQ7P:X66:VDM@4Pb7AZ.#c21^T(g[NHS=FeFO+VaZB[(W5H,TaC
5RLIMFPW>dT#49E=,bJ2cPZdVg9R[9[+E=,^-L7[4,7UaBY#K:@:KOEMEZ;#eD;=
X:=KB-9<9#W#R?;4X]N;++5^5P=3:QT5G=TOH.RE+Tf+K67XI8\6LJb:a<9[AfTB
bFAPEbH9N85L1;JQ3_&KfOc]PS:D2\PXRPSNTFB6@YBdLEOA,8B?/B_>;)bdS.2+
]^PeAfA44O3/fef_64a.=HCL(Q<05UIRgZDW[b)[CNTV=<-Pe]=.&51ED3PeAWYD
^g1dM<B.@]^8UI66c.<1-VGX92,;GQ4VA.C7&2ZX\PLFPe2][U&<97A6O/^\f)RW
g4VaM=eK;>Q4#A-POVN)cIVJ]F\#S5Qa&M=ER:>#02^g;5bZW/<Y^+0EcS?LB1e(
,UPQb/M[,:14&PJC5/]^VR+ge1/^V?4HfZK4(7G-d>QD0Nb+,5VLIML5SRafHAVN
3VD]I/=U\KgE5aT3gcA7Q?(a2VLAeg&94YWDMPf@&CIHNO[6FN+c8/;eD9[Ma8&V
cG=PeSP)d^L5H-g0\I+F+M(J?00^69I,>eA96/Y00TR&]B^X)30UY5YTFZPT5MJ:
D+^G2+CCU+C,-#5=HNTQKZ(J<7X)V03M=,I<JJ=:(gK_NB.A\SE<a,/WJO&@7D(C
MQOb/<b.Y]gYZ+OEA+eUSO;[OdNTEJ[;4/3^Mf[T-JN4;Ygg?[B3aHe;BK(I)]Q4
PQ;cVVQ:KePYDOe#.N0Q^=)0b996N0C\(]AGKYJeF/XcfM74I2TP:8UB)SQ9+QVa
).c.a6:)M#QJ&U_E@77UN]FZ7>V]7,4@U]We]U)-L1J4?+EW@R-^;6BNgEY5?YW6
//_1/:))JOb1aIe[:Q@#H[GKM=&>)]fQ_5DB_e9>_dJC5HdFgD10Z.5=CZL-+/W3
4KZ]9V&,6S]&6a#2Z>P_O^3BHJL[c_V>#E+42DUV21c4egEFc4;JK[DRaeScB\BX
JEG1?Re]e]V8Q[W7eOU<F5Of,Me1V9Qf&BARS^1?6T:ca&gUSb.>Rg.58e4Ya@=^
.0<F0XdLA;M),?L)T4#d#4gTG[>3B-f;6IG\:RM[1/<PMc+a0aZgV;]NL;)3F1V,
_Z(\\0<XW(Qd<E@-K31;QNF&8ZF-7ASGL]Cede/8aKHG3@YaR5UedZQ-MIKf(D<8
I@0Q>VJ0/N-:#7EQP>XE#Y(UN#HfHEUXMAc@E2dR2:<Q##;N]&T785]WK5gRgKe.
QN?2QKcD5VdILSa#(e9E&O;<f&K+ZPc1J?Rc@ef9/fbK=0KbX#AS#8N,64Y,US3G
BRLgW5QY6WJ./R@@T;H[BT>4W[+9&faA/,JESYO=CJ;#M)dcY@Wa;=IYV_MOdfPS
D.H[b,?8^55SU#/CbPc2UgJNRN1MAXeRea70H;Mb>,;7+=7R^OE<+#IZ\3,3Zb62
REH<=20VODf0YB1bFT/Ob4->[N\.--YS^TB;?]P8NW>@96HO(A4_^2@/C@+B)XO@
PQ2,N(0B(/UDU.DZH:9H6E,MR,9PZ-9WVEB2F4b6JSfg-W.LZ1J1d-a]?II>U\Wb
G2T1UO6YN+)J1G=58KJ1A+=^<-Z11E.@f07;.7=QSFb2@L:)H&/aa\JAE@2+4d&R
ZKFQA&8M8:>9Y1^J-7N]M,^JI2,&G19>SL8=H\23:DK7>SVRfG_a?OW26;M&MUK8
bEQ.;W1HQWFRY[V]T8Y0G:MbD0)?L/CSHPU_g_OP(#>9OHA53QaETCX/FU9\[DG&
2AAV>FUb:3>ZH_F]bg,CTS9-N4e/,Wf6a:ARTbA3,#(g9WK\S,3f@.[_[.]bcT99
B_T[O/EXcf6:;_ZSX2>JF/>DPAHU_QZ/[^8+&UP1?2X.7[G<e=D=:0Pgc3_0+/5G
JVYI8Z[a)7g^aeX(/>>F@\?)Wf_YYbWO=?1Q12J]1[AHZFPOJ?C;ATC+60(FO<XM
YG9(J,SW+M>MF\G;ZF9N655Q:(Z]]HS.,.;GX;fUR&1/,ZST6XCA)Y@eL4(P\e,Y
R3+EBBCdfK8c&J@0SW32Z.T>>.J97Q=&.\7/=8^Y9GD)]e)2F1>3MPZD;=[HJ6;Q
gL>9+)R^4[AM1b])UP#/8H@a/,AW3L+44UIVC#e+fXY[KO==3eXfGT#Nf^Md0XC2
TWNM2][EBCag4U.ZJ6:JO>N@aJ>15E+20[5[g,MG;[=VbT)_d/c&;[D2]/7:cCT]
g#fNYfcLKeX:HSf@?[F-CWb)8F8-+NJ)Y[-e85:V>+65e.G^QbU#4c-IT+PfK@d4
G\9CB\ME;1[M/c<#P4DI)(5[d8NUCQ5P->A35#V:Q(0XT&-<.X@+UW6b)9=LBG&\
Ac[RbY8NdTf8)C,HdTc]a9QK;cg,(@[^9eRMJACJ.)TeYFBdcgUSS0\6Q<9UP[)M
U2^6;dE/fTF7)#G63(/M4Z^M+I3A^K\17QU3/dTDN:a),MIIRZO/U]fad:]JAcOW
IS4/LT;<IFDZR^g)0:?7&>]U,R1C[\WgdfWfDF+7WS&H7b[S#U<d&>N_YDbTZ)c4
(W7GX.^A,:R<21>?,AIZ7HD,8K2VT9_#gY\M>c+);/&O:-Vb3:0EJWM^a=S[<4>\
_MDU>PfM?GXGCO3?O8bQbH&?7]/&P2=^P?H#SXKIbJN3R-+0E(FIU<5<??0=&GN/
@KYW[.^Xa+F5W6YU-Q\<abQH-c74<+2MLHSRafZ6TaL+<LN7U<9L1fR?f17^^\.-
5[7J];?1PZJPaAWf;(e0cRQ=7&EC^XI]Ld^=IB\.c9PTcE.(-(TK9KgB+A[<eNY?
\0-WbDD+EDCE([^3cLdFHSMCO6T@>CP7MEJe,&TSDC>STN7A/bZ^S1bIV[39<aH(
-WW^,a4&P2D_aLOWH5,+F5OD]-KH3+K0L4&?&?NAbc@ZU#2Kb#T<\AS.XE^fA/8W
T=P>DIP/]e+KAE=PC5?RCca)1N)C(/RD:+A9]JJ3/UW06W0:+4Q[.P+Hb./GaS^a
[(#<VE)(N2.UO&TR3K:#aIa#KOa?VVKbJP)HWd@)f2c_a[2P[b5VTVVLSK#@F<E1
UO),MQK6dVeR8)FgD@SW.<fQH5f0<7RNfCJG^d-[gS2+8CWZ/QBTO?P\9GJ^;cU=
&M6A6ZeVd-3W_T1d^eD_R:()/[I(7)NAW28W<OSa;\0.2M0PI?H).ILaI>+:VFX4
@Y+6,0fY0A;YFECU0-bS]J(J[D<O]OE/cfF,U@D)E=#&0;\]DC,_6=g#JRDL/,O4
4FfGH&;TE<6-:<41D39A<=??26<6Wb(^d.dX<J_4//,2;ZCJ7Md3gX6(8D-2/DR_
3R]2dR&M4:6fM3GB<VLTPEQS1;)HPgJ2F5b]gVNK]gTU@R57?^J2K:,M;]M5,VUd
EEH.b;4(Y8<Hg+&@4SF=6e>5-DELC]>-Td8NYR&A3:/Q;<:F7e1C4)L#e(9(U+F]
SfLG/DHTYT.?d[93gX;(>T1ZH[e8ZF1XMbF-3L-(f<&S,,:f12:9;^IRXC1&ILE7
GR..Y#IO4<IACDJT+MGV[(2IQd5e-[+@))0L#AN=34EIG_0@g3DP4Za,V>N:]U4Z
Y=;6GQ;MAgMI,JId2R.VDLG:9_FJFO>(FR1RPZ3H5AbfW^HV4TQKS3\:.eD(M8J;
280d/-d?&+?#HBG)54eRR1;P)K@9g3/dT#S^b;f>T?>7^OD<9\TLW/HP3C=O9S=&
:0MQ=/M9VOZNXa7#^O@C-6QQDYU?\c=4>YY8MN6aY#U2,4-Hc^=9ea3J24/@Ha3_
cLJ0_bLZ45F4B_(g7<-(U+g#^[L1DII/U7X4#+=f19JeA9R3&ON)ZU0EcOIf9B+L
Dd4)DAC2=#&cDLW;>8?D6aQ(S>GLcb8VLLHBNE=PJE+-6@D(X\;&_GW^?B379T2S
cFY)<5MXf-RYNT_6KKGR_W;I_).Y\/>+fK,V=5+#_:^5c)DFbYCGNA,6KMf,\UBE
Cdd,3C@g&aH_dAIMbN)<5&Q#UGHDPSA;+D1<(N1F=H=a\EGK..YUX0aT[E?R>]<0
?aZ)AM(aH=\):D@L=Y[:U_Od2QU[^1[e])T41BaZgeZa,K;4OX.:PISJ:7DEeIU7
MbceI;Z.2V9f:E0a4IfbU)U7ec;bT)R\&RE5WWT&G1RbB5H05,X)+XcI=F09Y_>\
.9V59YWge2.SgLFOCVg#7#GX[S##aUH>3V[GaTY-&8)Za\@9^HQVD(R5CVfG,;B0
S8Ug?WR&F.fUE7HG=#gBZ1Tf=2UB\MJUcS]-M_504dX6U.916ZQ#_L7,/6,=NDZ4
0-1>FHHK5TKeBdVU)A-JUP@](C?]#2Lb./U:PKQ?<KI7@D[#e=SYRT;9U?=U5eJ@
c;dI\;>TH&GfW_O@Wc0\Y-H[-3Tg2eEcDeF8S=](#ZEA;fZY#>.XOVZJ>N&BY26>
-d[8+]B=GFC0\2PUdc)10/=\Vg^+43a<BD#=RA2M5?R&KJSf]\H4_60XDQ2WC(W+
_9FVfDbRCWgBN)#ebT.OPHe:QB#Q;CJ_e3WH5MLBS=Df8L:88dWe6&>JTFK6H#1G
><6:K-6FJRX12-M)R?O9BYIEH#=T\86dbggH1=5dg?d6,_T=@Q<#T>>6J8T+QfZ7
\PaA+R=)/RPR7IZX&.S?BbS;)Afa2)6I8OZ,YbSZJ]F@d5=CB3O&.TC95g&ZD<-f
Y]0MF4Ea_[IUZfLA=P-ZX3SI<Q.eXH\;#e_=@daS:6J)E[XO<.WN;I1H-)LK[FCG
.((]?Vg,K.(>U&8CB+9Wb1(B5C=KLGKO3U5(8XTQ/DH.@RWM/[GbD?eBCMPKL#O1
Oe^SB]EM-A+XfDU_HI5fL5N+M(5=_89ZZC[LY\,(6DF)-HD-ZU0-ed5\-ZYK56E<
:RWfT?Z^,?F:TN,.-RgAFG=7c?>J@8=ZA?_X/PQ9MR>[dJaJ,b@UfFA+MY=]B-fP
)&5e4IR<\IT+1=8NQ+D::CFQ<L42-&&I<./XC+&65(L._LHWGg,;egG,KDe4=JPb
K/AH(aI=T9QZ92A1?DXUBIR[b8@#QQDZK+F]28X)[7@M7Y2[gE<P]]CAc5&^L:CT
UVUVUZaNT\5GE.6ML?YBC;_(FB5?K6QXXQ/[bH]4/:=]\&ZZL(D@O<.=,XA/78_I
]\7bUA5K#_,&DJ1TPNJ_O2f5Xa?HKZW6<])?[VC#H>?8^HETf[E++J1[M5)B74\@
CO9)R&,NX>L\AYNWFZd+WEXD?S5XD9#;^bJbD<AZW@P\=deQ,YBbgZ<K(IaYG[\;
04_GQZg33S]\]+\/-QK>#-^C@1)TY?<2BQAg<Z]-1K7R;8JGcb\G;?(HTQPC8-R9
[9XB7S,ZL29RA.(4MBOc-NH7[ReAKIG\bJd2XF;GE.Y-T[IX?M1]I.Q<JO9GLYe)
/C]cT,<\_CC_^c(;c;IDYZ=;JXH2Eb01(.P@7FGBL?DGaSOXcL3bQ@KQ.VPMK)+(
]459[YeMPG5>TO.d;/HORTE&<+UKg/K+OY?VCN;HWL]VFJT_[8MMVO7Ec:V[a_4=
/.)\T9X<Z7G+1.OZF5E4C1F4f;dIKK29R;AM99[;Ng0BcdOT(6L^=5E.@(XS6)OJ
X39)1F&Cf#MILI#PVCF@^FadWU_]CL?KX:K2D=&D5e9K/C/]RXf1PVH956032)LG
Zf3H@^+F(N?_MA;Y[.Q>=UTES)SHeGa7)TXg9NdW?<eH4M&=@9G_+ZVXGG1H[H91
T\I<(-G^1@A5:I84a.O#C8/C.bHb?0b6-UO;:I6Kg2GTL^?C3E]RYGAc8Pe6KNK;
T\TRTU6CXf#N0ACR[EL?8E)Wc.JU42=E+gfJ;<&T-OK@Q>ca<O(AEE0W6KO(aE)Y
_g+S,U6E<J(HJ/eYN?cE0FP.UcVRRf@eN_U/:7/EC]\45[=NfE;C<LKfdG,HPf4a
YVeO=7KY?e\9Q[8FL[4@e[:DE-[U=XKOXYSZQN^3C/0<^@>_ed63CUfS\f5T+6QT
5g<\DWHP7^YOQKFU.^Rb<J#UA^PD#QL#O]#<^5IT&b:Ib+9M<+K3a6HMb/]]3<2g
.4T9cb()#<?90S@(KcZZ^93S>VTd6dPMT&J>(4@^XB;KEd7YAIE9TFB6cR0&&I#d
Y@^b>(2O41KY,YDa+=@eG#50>fT483OA&]^^b/Y2e1/EgW[(J=JB=Fe+/B#YW.EY
eTKI;.5-HD,D3Qf2.Db()6P7S3&0eHcEV,f5eKD<@VT0MXfWFcD5g>[2RQ9;dG;/
HZTZCES.CPZ2[3AMEN@QZ/[J:5FF]A/RYdQ-YAFN].cN?GR^_OBe3BTO\d[M]KQL
Rc&[\6.@(BKLCMX8/I3c9Y\M,S/<20=;.6&B:C;50eEGVS,F]ARNJK4_J=^g5A8M
BaaS59KT(e[N?bG[[?UVaEOFC<KJ2;-G\9._^[B\+(IfTJ[CWXEB;&b1X68BJT8R
#\aNWS;FK47O0+4Ng.I]GeR&_]1G0e+d1d_gHDD])-QBf+,01>Y)](:+O/5-IeM-
=H.#Q8UbQ-=IRg??9T==VacQ>1fTP8MA+J6Z>TcX-MQE:++YG5GMX,UCJ8FO#WHf
HK)_c8TC22<2^dN@?eA=DQcG1X3/5e-)\/:VTL2;P(LTU68dE,C]:c)GYEc75D#?
da.T3P\OaeAPM]RdCL18JRb21+MG3DXP\Zd[)MO0X2aa&OHDe:63=JW7f_(^7+5R
^)C6)Y+bM&>@a#)X1=7c&J#]J,5Jf45QK83JFPc<]7SKR4R<7deb.B0PQA]Od1FK
J\GcU-K0=a\T2I@\-B,G[MUgA3MSQ1a,J1YHCOE5>25K9^e<0cb:#+Z8U1VHN00=
P+d0\F>2aRN)+[,Ze[5MbQRFN>eYXgR9d,JQLSY&8ID#GIJX^T[O2ACdL\N3K[LG
LB_U5^2L.UC17GI_QWQD<IIC;fW+80HM?8/7[BaPM#Z@]);gM&EdL^a?EEF?=E<:
ggDW-S+2CB7?eZ^&?I7/5f=)F8^1#6_\ZQ-X5R&=>T?Y-2RQ8A8GKK+?NbM\;Z^a
;(eM^AfFO#2d/TZdGbcXX_=XD38<<U]:g8ART^<VCdM9RF[9-=(9FR]d;X^D55d]
+(I;Q=3966JP&DO:Rf_8KQI2Ba]V-G#=ZUTDWJ2.>E;S@X8Y[7KH\A(?L].<)3G5
8VR7>M]7TbS)bI]9RF0Z_J)G+[KHMN):W4=TQG_gSNGH[5Y.V\@HHRb84f6H@>]K
&#7,7#E?bSF(A1\PC#<g,0Ha.I7P:+2.3A^V9UTNA<>4=027F+QPU.\VN:HT@@+?
]<?Z&WRD4<_-IZP>9^GZGVM3W77WY:Je(<X#N8&WD+2Z@EDOPdfUI:=8Y?9L4O?a
;SWQ2Wc_d0ANY+E]JWb&=,fBK^]Qe.O.5NY+0@H76&.>#+48de\03Pa38O0]/FB/
Eg:3_GIf70fHUL@&-f1SeK5]Q>Wc@+3>.WS@LDUdSN=]__A)b/3eS)_F>[\4Q;ML
L/Q/L\)(QdYeK6QZ;:(_I=3(8WID&dcS[/>L<f)GID/V07OP_Q+3R]):Cd&_R/?1
DF-?Q_NSP<e3/cOb.3^a&YcM=c;Yd-,:<^25:8(,PGDJQLE7[9J&e2LZ.)F3FO@2
82I=BD0gF63AZ:<.K=-6c+0c6ZY1N-=;Tc,[A:]e(UIM\e638Pc3<[+18R3<?^6S
AeHaBS^>TYQHeEQU,9(H377B6673I)B@-G8;;8eebGGfRI@/4)E)7>[8@dZc]Z[G
?JLW45KQ3UZ57228^M=7V8W[IBX>@d_UIc0;G,&DVTY92TX-N1W5J&2Gc[4#2/gI
;2XW7E9aTCeMT&Z@YJK#YVD;D9dg^Q=c;0a][<EbLN_.A?_J-abafKW?@-P8Bdc&
&&HNA2SW&J)BZO/4]>Uag8#d]a^E\E8[K[;-DC=KAdDZ-6+5HA+b[aeWbSBgXBR_
ETVY:^E@daOC@XD2Q@Lge,[bGSAC4XJ43#C,#DK,4HR1AZd]+?N4/EeK049T:b>7
-C8^UDCfF;2YXKR=cc]cL^HV(O>LB;2R;6?M2Y)SJ@<]\LG)aUDQ=RV:XQ:;bJ@6
XH4GgdfJegHCS5e=G@/H(ebPF<1GAZ);(KMERcDg3I<J617<5f&M7)9a@]+.;]=@
Q[3S)?D^5PF+KVSIEF.IQ[=O(PQG?I&.B#[LVBI(6b[.\[ab#QK9P9=F^\@S5C?8
K/M;c:Sc1H;Lg7bA;]P:L9[T:e@=fY?L^KaMA_NJ2,7U)cOH1:+5LJ[1(BO.X^P=
V;C+Q4L>/6\]T[X3DN5A:YA7911NgORM#^+b4CJfA&;1(,2B:8IG=QIWDJV?56eO
7XCS&CZ4Q:BD0d@WgLG4-[@EA,ADX79P/0f0?9[;WVb>46&7]e[O&(1gFgQ6_5Z1
Y<\Za(IaT6(7K)S+ALJ:3eE)/W1T,PRReY:/Kd7Ue\,@2QK-?QJ>->?-,[SW@V0M
#GSUTM>T25g00C;J3[Me?=WQMQBZLTGEBV^&N]e7@\]4]7a5f=_geMG&Z_26FS,7
bZ//Bc#)b?QGg\:7a;?QbMGe>8I<)AI<Uc0E>8]04B];UE<;D>3g)S+FLL&6[<Oc
c[YS(^8:CD)LV7gZd:,.9OF:?f:7Y3+ZV;XL737:\50F;SRR/B23cP>6001#3UBg
>DadLe8988e3CM/-f;68+6+1@J=+RDN6MGWd7gWE/f(3._-V:8b9,.MZ;4e6)a/:
b4,W^_Q>Ba017<\XRA&S^AbK(5GS./d:[beFC<7YQO]#4A,TZK.;QBB\)TX@D_1R
8@WP00KO;?._(eNcW3JSV@JT3Y.cJ00SZN/&Z1b=9/HOS(9+S__d/R/30DZ(>?R2
fH@E2/WJ])QH@Qe0SP^,&]K[dcZRC13KD-H3KHOKO1JPV>,4_;Cc):aS_EKT<2UO
<?.7UD]BV+-&(C/U.:(<=L(PQP9(@]Z.>5G#F,J3H8\gQ0BZ[Eca#Y;[DJ\VJ-@V
;=O(M>.dgd^G(Z\(aDUfeO\_ULKg<g\90Zc^[1_VSa)FNW=;ZAe/)e>L35BF4]\=
gNUaA^JD6NSX<8C=]OQ;Z5KKEMd0?JB-VF_g<+@+.-FGN_K#5_bD[dSL]W8QVF>E
18]I9J>e=fIF==8Q3=2FP?G1J5gQ,ZF:4<[f,66ASYdNB3_9BJd48-65?3,#>PC]
8]8b:S8K-DP;eU&/?[4^-?V5VeGGTKJXRD9ZAR866DdbU9OHEDU).[DQU].I__3/
)TK2AZRW&#]BFHNf;#/YB[:,_I5\Oe_>:9bcIV8/bMWTTW<f6(E]REgIXS#LGb=)
[O&X1(NHf.F1V31IJY#W+Nb^MQdC;EEUAHX>=:#V9C@)/O_:T20a,M=+PdP/2Q,5
d[:&Kf.ce6B?L9J1LWCKW40AZWW=2.;+dBR>9\WbfI9+I1+E<<F8-f&3.>?d9\+>
YOb,_HFR6/#9#S/\X#58-\J8P^N:H0F:2^6O@B?ZUe3Ke\cRTEU1G[1<(#dV,EfE
PRC>EP,7J05E\_3X2,.Be=/@gN&H87cT=I;CW<Y)5D6A[M\He4:IfOS_6=1&WBS_
[YUbPd>S5c@e.G3CQS&:eC,c,P=ed/16^^6POcQeJf91IA1[O14_ZP5f)O;.-22/
fLWQ84E^:4089(cP1V-Xe3Y4T4LbRLRU(^X?PWfMe-))+W.4,-;?)50cBRUHLKEE
^5:RQFFJAR6-+&:I=A9e&DPSF7M??G1#3LM(K(&W+F^.^MP5?aF0G(,U@UKR.+9/
^,99bU@4OZc6Ke&S]C#1c11?<XC&BV9#W=Y=[+RW#J;@XbHf1_eFB(F0Qc<^0AZ=
cQAP(MS.gGPOg&\#X0&)RVLS^cQ@0NG6ZK7P124aPC:0c8M)bT1)0Q#6960#8M1M
#+GTI=gM(<f>WVQCgA.ISa<.]YDa[0K)M&-0agfZ3aQA@>TRASW@RSYdASOJ3O)G
.fLe?M34QY/5A^Se9149bJ5HQ=fdQX@H8B>cd_^M#3<S(cR<e(RU3L.-]c>G)TWQ
H_@JQRJ\V?[=MRX3ZP409I?F7-P<G0b:K?SD:ELL1/[f2M56=5X(E154dJ\e2KCT
Mfe&L,U4(1A.EX_cTWg]ZZ@:=FXffg?+Fe=]/?ORT+>QFQc(SFC_U3G70M4F,2<A
RMJ#63/8_1@06f.5-&3G(=7?Q)448]:[VWDG3+0dUJ>\NZL-)IKRSB,OY#I=1=HO
P2(:^JJaRMI]=@CWN^GZdA#NVK9+6>(9;,-NKCd(08&ERC]JOC?HFV3O]L?ZYHIL
a6,Z,V[<0-3=K\R0M9/Z]aB.H>Ag_g#g=0Y,f9FPC]ANQI,?]+Eg8V\[e@aTN:WO
+QOY1fT0fE]DPGO))-G2^)<+U]g@cZFSN0H@UYC^?MBdZPZW?8.();8Xcb<GZ86,
OLe;V/?()N)G_6gFb&f@:BWeO:[X/J>N0(VT_>cIMOK2;55DQ-F1f43M,@[V;B2C
RH619<IX07#N@>72Y\IHKJaVOIHX1_=F&TVJ03^0W@W7/IF1UO2>RIAe[AEe[U(.
[.15V=>bSY#TJU80g@aJBNUW.:08H2+5cC6Ge#K0[&;KTJ]=7@2]eZaQH(NMP<[c
S7b^L-EHOTSZ,&f[M>X)Qb^00CSHX2dYD_OP=E@H8Cc2-Z5IEWG/^;&2BaeY\5QJ
V?+X^J5-WI<6@e3&7CZc/TRSWfFK5XbCK@#QY8_g>]XNW9a)0c@SR(7[^TH_/6._
?3XcMaHH#1.M59B8^14LZ2[=HQbBQ8(TG2O>,+B]c2d@G4YR@;G[-4(OSK,GZ)PK
QZ>bE&e>01B_1aUHc0NP(OODO7TFQ<JgB>@Z@81b_@A5Z8;aRQWJME/_@88(5(a>
cW[?1Y0@TeRY0_:L4QV-P7D(B;M:9a7=O-/VK1.bL/OF,);=cM91YJL8(AC0-d:B
M1BK7Lg6e@c]FCc<X3Z)?A+124&Y5YTNB^882Tg3<V>6.>-(2LQ2\8>-C6Z7gJOI
8Vcb2T-8K+Fd_fV#6AMfN+6^.)-IbBE<]UHI9,2-6U/I2fa78^6P9SbQ8DWR41-<
6Y]N?VJgB@5E^=ITENB?FT0O\gM9-]L@QfJ+cH-)=0=DNNgS@Y2?]K4aL,U>(dAP
g?=JSH3:CZ)RM(0,=<Ib1OS;(URH-NU>M,,.041a7M/-C5S]HO<OHDK,@d;_5G0F
,g<D?e)/-L9QZ)T0M^X@Q[RB9KIgfP]#QQQS8UXZ(6Z@F:G5EK0_J0126(&4Y:Q/
;^?X^agQ21VN9.Y]E#/a0fgL0\G[4O>J?Z[DW:E05O0-^U9VA5Bg5I\b,9.2(#KO
Z2WYKELA+<]N2YS9K@NY<6SHFZYN8V:Ob0:449,A4:K0OULa,^9L#V-GNH:QM.,R
V.0a3X2SZ[6f0?A6QBC2d=P4-?-(0\9MFfe>^?)VB<3_Tgb0QQT/AU\6eC<UXFAW
VT>gN-4,eK.;W\P=YcgV945XHO;A59HV01/)ebLA3f4,N9UBRb<?QbbNa2:I#(4H
^<<SK2D.Ec/B\KK2(Q&-(H[4)YX34_8d,BW^.]TAF:9;AfDdY04JLM_OSMBEccdB
:/.<@2<)3+_)MBD5I8dMQ-NN-4_F-+(+0fA6[?3Me\5.U[QJ260dIMXLV\J@S/-O
FIcC5<,)BIMX[@(3#_/2<N#?8Ub]>G1SV8b2Lf1EQ@^@a?S=O&N_0&?C+DW3eX7a
agOG,=T3)&H);?/>LEFBF^=4=,)2]Jd_GG(>KAN?:fbJY,Ma@c/B5J91g26BF_Ud
K6QeYZf8.-@AX>c70Ja-\6_BeZ&ae^aJc<^13_G1_ZB9<Ua./_?BRY\cX27Yg5Jg
;@88dX4MFXa&XPcc6b/g]]>^9;AA9^D_WQ/?;>>GGH9J@Z<QTfMQ8,g+6(@]6YXF
6H#YARJGbL.)I(_DaAcG3(+19W7QS_NP7fF],/=LTeI)4+T1[&=IX6SA:a?[b3/=
V2A22GD.I+?A-DX3D5DGPOW/K\G:Z6POdC<9Cg7c6GA>K>;3DPVe2BK@GJ.AN;\;
@^EJBCb9H0PEFE8.cX.3[3cRa&AL9KAP/)PP)XAdX9B-R\MS5ae2@[7^\I=dST=W
5gF]S5Kg,16KaSA+?J(aG=addd-9]NWJP^ZQ8W/bO<aRbU[U;SLW=+F.)1O/QE2G
;b)(<&5+Je&^JbLWV@WaPQ97<Z1U?,_6CY-bW#-?^IX,_:UDc\7&;a,&B:SgFW,+
&)X59=Ng4:8Ne8?TF@Ne#,98D#0Y)/=F_QW2LcFgT?;#7)5,:5D:.IN2(abb>U0f
3bbG9\4M>a^3)XY&LJBGI.P:BH=dE\S5P)3(S1(H:TZ490JMKL4P-XOA[KDKI9=5
1b@CPFg6=a:dNaX]&\\)9^4b\<@F1eCRA4U,=YQW.1]2L.Fb>Fb>BCO(N#8QUA_I
:JG)UV2)/(c9B.Ge\f7V(N<0[Z.=+@K,;ca]gFSbDW9U8eV0J\ddAF;Y0C)0C-M<
E5B=V,>=8+/0(I+;07EE9FaR\=&4UL7R_C4>):P.IRFEcW&&BON7:W9]7H[c>5U9
Ggfa_UI,e<HQN.3+B\#2;eX7WTP(8dGgO_cL;;M[6-_[fI>gGHcXWb&4X?/HQ0<I
7/N7G<f:@><I5BQ#\RYAeX7.5fX)&H]/)C9D,TLbc-SE>:8JTC596JRH=-c?^bWN
JV<0edL/^c=D@[\K?<RX,CXRa8X1Ad92T(RXRAM6S-R]J41.(ZMQWaa^,_#:UAIK
YHASO:UH<04W:b6S;=Q.K)aG/]E2Q4>T8_+H3[TDM]EDf.8c?NLCHf13Sd:Ied.0
J];CZe?C1]GF_<HR0SB:L<MK@)I1G-;-N2FIa(2WE_F8#A@b)49bKL&dSOBIIC0L
XZ-@U^?S7I@B(c34FM,-AdN:VP6cc+eaQW69D3Y)7O?TbfdRA9NYR1AR.]2(bb8J
B(X^IND/5P+VbMP)E]3d&8O21gR-AJ?149eV5PKTAAM=CBF@L()=/W^/e6cXXKIJ
Y;7E[X1E+,+6]eSFZQA#M#-1&T5^(1MQ4[a1KPIY:\Y5g(D^&&eA1_2L9Va./>X[
e&gd&Rc8]IKCa[:42^;,_;8,2I#-:IH3@2C(+91W#g::C/(6(Iea6WOfX_P.b_\Q
Oa+M([9aCH&_X?GP#93_OGWB2KNR:Z(S+#GT1^IF)W-X?Q\;5AF-bUE?=MQ/BBWR
[R&>BZAdSSACK+DY8a77=K43(Y3\gKbD>7bbX\>8c3N=/TG_EU<FU/KCMO7U(P/4
YJ0PDc,7R9O;TWa/8NI_.WQc([?>?[0]1+8C2f:\gR.L,4&Od3LH#-=g:OHR)E=9
&@PP8JXfZ1-g\?ggBDUZWUF_2#SWTZ@/S/;CXPS;S\dfNa3#S3d7WX,2dK/0a>#9
/&C++0>I-H-gQ\)gFX@+.f5.H._VdRgPT[;ggMV(#<0KJ_-<QWFC#+7OWJMK;aE/
L\G&E1/d3eN#03<ABENE4b0]d4MdHHR9-=0J?(]_#Y^eICS9QQ&B0M/@A+dGS4C/
-GZF)M[&0Ib0(bI[CLSZK6Y&cLNP=/^YJ0Z[dH]F.Mga,U[(+g^eB.e\XJVe2#cf
34,d5.[D,,_LH&6db3:<[_OY7G:IK:f5V1W#/a?U)<SNR+ceP#65GeK/352Z[Q<V
:g==aEfBV00Y+ff4FI@H+WTTdTS1c:Z89<#4PZ<8_^VY-+0d?+3+WUR;>7a_+8R^
fgg](U2\BLN]+<+Y&>9WU&ZWNYVSa7>A>^:.5;?<=4g9bb)<CGE0c)R>0VKBXI(=
M/T>=2fL/X,Ma[:(3T5Ma4bJ,0CLY/XC4Z#]U>R-g1Q9M91eN6HK)\?1X>X?ZfZT
#_##.Y+/NTHS-)C,XE3P9,b3=X/66XZVWgZbB8_\a5RRP/WJX?HT(a/W3Hf@_b21
@CX7P4NKQ7/Z.ZEaQ)T=22PU=-C..3-0X,X_-aZB?]YDcgLP:P@@Gd[7X<9f=e=P
f#Gc0J)?0N+FE(UHL#?RS8K]@ED^4>b+6U>IR7=HfeBeaUd.^JAAPA>d9&ZQAcDM
B+,LB,#L2NG75/15+JLW_A7[DCK/#-aZAS4F#FEV13ScF-F+e,>L[7U9He=+.eK7
82#eP]O0P4-;+FYV&O.\XXPb7294N+bW0U]O:VH=)_WD;#Y&OMZ0.Cb2:N7c)F1-
_32NW=F(XCTJXIM))(<ed2F,1Jf=eSCX9:4VQUEI,a@V+JX[FgPK._6HV:g&?A#-
6?/DNbO@#5LL]Y>]089@c2c/?d708DbLSAVSQVL/.^Y3Mg052#Y6=B[7097-^b5S
E[V-)65F<)=M8+c4K3f>>[7LZJ>2\9>PJ4<5VZ_dCa<#N=H6&U,c<dI&LKO5e96#
/9])YUT?NP0U)13ac;9FBF>++3[Y03Ocg,JQg\Y[67#3.8.]F+fE\+Pb6>^d/0cS
ZSC&dAZK<dX>88[JV[eOE=_)+,##9)4B:dI/.=d4?NX85BEXgb),3dOYR:I.d/8Y
#B7[bC(]L#RHZ8dDR&XG,RL_BOXD9VTY[:L;?gWFYR3B4O[?VK]I]7&YfeDO_[E0
g:(\WB5JD/U(bM&>U5=A3D4>Zb20I[-/DgYaOD;)+NW<9KQ&feb_#f3.(XAX6<@)
CH/R0YYZ;\.;U/WKa.5AZ&KF&GU7RF8FBP/H3SES<Of[5gLV=/LQO.(&b?.EC[g>
L/X(B8/dNI7YggI8?YA&X7Yc,@^6P0ABJTg1/E-:.L2<7S-0\gJ5e5aQeSHQ#89_
Z\M=;g.41CX(//Je_J7d+]f?C6OVeE^2>2UJO:^g00FQ\J=4EBg.ZP55U6=fSD4=
5dSQ3A44-gX-67U;ZWaCO?f,>5f\ZOPNZ=b6/P7;H=:IE)>KeC/I+U]2f;]H6P;L
IN=9EE8=/7(&g@>b\5S]?7LK=-3YAMA=?#TWWdV^42.^WKTM^UZ0UCA,YD[[g8;J
ZbOcBbIH.W3@cc6dRM+AO3)=C_,YdW7):95ca#0A\?L/ZNATa<YK-8#YVL&Z?=8f
,B2ZOeC1>))[WG9a+,,8C(#M5ENB&d^T.eeK(O:E712I+<Z<YbJ&=R75@0DAS;+d
+FgX3#D6S;/97-Bc76&1f5X/L,14Q^[I#c(R0WZ12>bY=Ae(G)112Nb)Hb\Te+I3
a^FV)3V/-<@EVfUX)?,S@;>P:(e1(efPA(IAa^WRQR^ILZSd1ON1.32DcJ_R_68]
1_ZHfUWJ-)\\0fDb7YXQPS7S)+P<(T/IK?6<E+f85IPUQ_O55\4F_L)#8U.PD;c3
CDUJTO^[LHe;Y8CGA&.YFd;fMN__:.Q-P<:+^,.EX]N9N_bI6OB1&.EH54DX].d9
#6f6+DOC>M^RBFB.&#Q?^I^BB)c?5+ZY)7g6P\gbNP_W0)I-KOF\8=E/;W9IQ/(Z
.dc=^SK:[X,/_-4,9<0F\^c6+4eZ52bX0UXDS)+=@7L/39/0P76P3gWY4V].>cga
Sc^BMF56eP?V1W4TRIM2,.<TDZ>GNI=4g63dRJ1XE10YJD/_KC5ERcE@@?R:#>N(
MF&4]#FDWcbgOH?<).dYT1&(WA:KJ(#F+SgIW.-Qa?]6)<DTgCH-K\_Ic&7PZH?#
fc<J8?a,,L#YO&<RY2\?b1gF5b@_#PW+USU^S5QGH1OO,ZaL&a\T&ZEM=dD_b_;O
C@PL[57>(CB]5e.-d^=ZXC<]c4e^ZXeIP8A5X@f)6dN@C8.<T.Q5^bXZ3<e;)B#L
bI)\G\eFGE\TM<6L<Y1-6?PI6)K<:^M1g/W6:G.=G4g=9SO?9JdU1+/\aK.MLeaL
+S@+dZ-Z&PP6@MA=d//cO#/c-4Q_572GgYH]Q7TJ^RXaYdD^FaVfNDG6@D[a0+Z4
9N[R:>OV5D/G>9WM/75O+E#BGe.VeGWR0MMU]S_W:^&+aSg]^9aFHc?a_eBN->:P
ML(Y[I#61N3?6[@(UE/16<_dQSU-B]bK[^4<,,;FU+3?^<;+1,^5V9;f8U44ZZAb
XY;H\?\\a&SbVRYcDKdd-@1D05DF7I-QO-MFCCN)PGB0/9L(F9HQg7FP5B[fA)L5
#MVV;Xg;?dIEFc34.5Hg__:NRIf3)2))=3U>-DZ1B>X#WJPcIe,#VfN(18NQ;U;c
HcQITHWSE</d8>5I[4_\aL.FIL=9;4N]C:7#,X.>.L3e7EY_W0A&XCKN2b:b:BeT
)f+CSK6BBWW^aV-]001BII2Q0KU@F4H]018;\.<DU[W378f>3GWOB^b^H-<ZOQ>:
A@FH=e>7dD8LXeQg62g;TBQC2<&Z+BddALFX/,@B7R8[7N50PBA>#?+4=3a#WT=7
/@b;AIRf4BM^:/gR_D4&NF5f789d7@HDKCASD/NN]bG.YX:^LJ7/)K0Kd:1F<HS[
Kc8NNO5d^L>W=+02:>g0\e7<((e5CC)6/0C;(a>W)d7LY^g09Q)I>.Y/+U3QBPQX
>eS?Z8NY#76d-C9UAA^_=K<+PA7;O\;?YcZ65^>V0O-f#P=+15.>L7&+TY\](CFF
-.gR6]FI1Rd2^E\XT3UZW2b?K(/8[V2R03-d&FI@T(d[LL\WN@(6H&bSM]6(Le]c
ZOd9Z?9aOWV:GbM,cAe(PQWGeY[Wf]9WQOc5:0>.eVVcQQ_\6N<CdaAdO10XJ,9&
;4N,#@&+H;&(/,^5ZCIV96BJHX6cF];,8PJQ?aXF9GUb8SI^7Qg^8_eF8,<[_Mf:
KbWYH+(GS(,1X=S6f-YX&Q;&e+=TXD<-/DSfggb@SWb>^5Xg#b2[6f@&KPKGL[M=
/^&YMUNb_feGW#3O6<7(U6g4.3=U7W@d<1OR>a?J>@=Pg:.Y/,C<,acgeJCDZ3QS
HQSC#5]Q<eU7;4<L]NMVL+:cAgL+6@&HW\Ye.R((HbKaO=<\.GADLd,c3G#cI#7#
9Z&A=LQI)X,YI+]eG_^b0OUFUZJgd\O^XBI,SGCKfK0,+EJ/^KWaP>777Ff.f)@a
[R1SLBI:ZR/)BFI4A_T+8HNU3bNfaX3AW2-CW:\P7Ecc3Ia3IF5,A-D8.KSQ3SR[
JJAgKbUWeD&E>TDA0V&Z:WB&&Gg04X+5HdS.3.#YQQ8Y##)N^,7<\A_[6&YLZB4W
1V)NYZDg;\,U7UX-J/-+J9B&8$
`endprotected
