//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
mh5cF1/DB2eG6hDExv7UnzNhnNq/x9NlO+EA07vZ2oZC0z6HKvLkblvUephOr6Zr
jq2LQxYRSMIJmZFEFL1Yl6j8vrxSQNm9bEBhljAHAsi19YHlHig38DgfvEa45KOf
Lcs7gfpze8gH5lwJVOS8FvoMCCMp3why9883yn0Zyx6bJs0ekm7tff3nApWlhAGa
D7b37NjJjdowzzmJGx+FhOD1rKk/OTavYFwpvCn2PzLdVc0FID1kEcD8xGKtqdg/
Dfk4Qr9ddQHJCHZ5jEymSWgqFhKPlRzYkD3HDq5Kuwx7G/Zh8lUB1PHdse9g/fWl
U8+TxCDJRjsd402pkqjSUw==
//pragma protect end_key_block
//pragma protect digest_block
wFt2EYn4QK+UXqZBJS9QA2IiPGY=
//pragma protect end_digest_block
//pragma protect data_block
BIx/PXje4GrVWuD2QDOpvuGvOU58Uj3pkT+D31yceWA7yLH+1HbmQv6ZK7zlG3zd
fF5UaOk/Ji/FGf5WhUYMGFwMIUGGp1Fg6Jdl1pIFTYB7sCFHBDboIZRsUHLVhqFT
wU2PQW9e/AgmD3uADAXEKw45ztzx1m/f9MsvpWeTKSJB819hhSv7WZ929DO/9vCW
YgNnqsrWUd737jMyEZYvOekCMwN7Se68pfJEBN/5sixLh9UZxRn7dgl57+Wnlqbs
mXAjvSNXsWS0e6vOmLpddxVhSOedKR5rnrmxDNZ7XABtTR9i4SJ7e2O0y3LuHs1J
s3uWEYV3kShF+Sz7NieNTg==
//pragma protect end_data_block
//pragma protect digest_block
SawKZhwavVIzGMRtLlYBHCVfqW4=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype.sv"
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
JvW9SbB7ReEp7ErydWgCTLsw22IUHvJYd7jjUgNEdwKgFzMCiYzeL11unm9fySb6
tUXhFacMI64MuoYa+TOhK6SsJqj/AQpOBRCu9kOlm7uaKvTj298x7P2loBUhP5V8
PlUKXFQKnwIX0CL/A1Jus5Ih3V2GoW1RnnxmdizMmFm/h/OziYjeHiZvCQcvmSFy
tRc4cBGhaAuhNZBWmq4ncGD/HfeQ4asaTvKIHb9yVKqPpgDss5X2goag0SAYWY8B
jZS+fk9KSQx8imqE5XeCAChDuGFUbCMgQNyvojBQPTruoPThxZZ1NrDrxcID10uo
p921rCMmb6+lvS+7ATRXVA==
//pragma protect end_key_block
//pragma protect digest_block
t9Ou1irc57bV4Z0bif3fQILFjos=
//pragma protect end_digest_block
//pragma protect data_block
TIh9IxH+iJU9/9M+q2wY2FLDqI3ug7egoefnOfRyQ1amfHhp3RfmwDORUVSKzA9H
VErCoMQNlyMX1Xa96mXvnzxMnqUohAy9066+rr15NuRkUhli+W6wmT6kwn8H2S8s
X0L1qiyPBNaT8bUG5w1mLca4vMQE9yLIxGg5sSCMnt0HldtHMynYur5LGMhKTyPI
I0I7qus7Wtg4MbH8BnABvMKKMhjVyqkUr4LllvA/VJU/bo1DGfXKPMbDCPVw0uuF
NhbcyRdX8S0OvT3xGtbeJMRMTxHhSIDab5jO2Q6ccb0jyrQN2aJ7OgE+QYNSZ7UR
/4ocYMJaq7tJr40HWFNK2hMncxQjAVCGEYwCke6VPEGh+ktZUsWN6SY1xHV4B3Fi
KPWLFq/tOQV12dA2zGXoFpm9BaPD6iX8JiJPmrpPCmJ64AxnkyUu5VvcTpHzljLS
w0Oi4osEXQT3a1ayNMI8rran5zcU/lpXNn64Wh6JBeO2We0JAut+PRbB8QP7vutm
43ffwRa8Cky6uXFcklo1LNKP+LpJhR6nMqOOpmmUtnsVbyaD20BE5FNaQmmKHciQ
LwCEG61J7UhwGbxXlsv55deDs322hB+Zpt3++nIFlbrCAX17FyHuwlGz2TAkg48/
tSKPEg/Rv8FSLOKlf9FQ5d9Xnnb4HI4pMR7pp0jMOL66O2unhi7K76EenI1cByd4
h3HSE0+bS/ICJEwKahbCD2B9F6L2OqF5iNBSJZqu7oj2e+Yhpa9PAAlU8u/YImNj
kOvZLG05BYInkaapgKaET5LAxuqmsWNCVpeDDHCI9FuQzTCcy5JOe4WTDspZNoWA
NCzky27wNPXSyrWfE9xibTHIK1J4m84SAv4zgV/byv8PxHuU9Feuc9Rz+8kKJUGe
2i5h0Ej/f9JhwwlSSgwdspxU5hPl1oRkELhd7ysgiExgxmH0SkCZyYlpSG7De4W8
rtiz8yt8WCLI6A9wuq91w4pMQmfIo2i/1pwi2HLFBCfI7FPrSNrm/7HXv8lZhwql
TsCo56gH5GmMYzYfD0m/R0ZBVFKbVbVJEgVZwQ1XtJoR649DN1/jnnECMCbEjUun
ec4mwPbcRJtZujG0vgngVz4vjSxR1taEyaoL5w4HyJN6yfadMHD56+y8QqTXzEes
IQXNq6R1J6rX9qVaEeHwO4lWpo0NpRLEKaK7f7J2r5LYu1ne4oCkFh5nZBkuSf5T
E6B+XWXJ/j3Ded+E9O0FqwwCGhUPuHLu2zsa7VzJOfKSAPAkAyJgc1Dgb+lKh7a7
OcX1gT2nWOZWe+VLrgDd1K9iW0HPJzlSo6v1Uqd9js5rlehA8vGrQ5aL+aGlxYj+
VHV8DNT4AV4iQrteQPpAtdz8g0Ezz+7mkSh/Bn3inGmzmOKeF82sFiLC5905+tX0
BM9e/dUS/xl+2w423B/4DPa3LYjrHheoHcrlRsyfNvWeiQCz3Hrv5SdCr4ub0Z92
DiujeImf2Y6J7kDs4bvAYvaZ5+Z2VzUs3GiFKcJAYnxy/FdnaQDNVQEa3e1ETmHO
Xflsgx2LovGy6+QN5fipRJ4prxOp2Elbcnp+iIzcq5kS0r1vYvyDDGdJeNitDyLS
9Z3M1/QFVt6lAxA6NmcTqLoKC4HrtCRMZ/EvDqTPWAnLNiS7gqfGubGUdo8R/7uz
mkP0zSWWhhIEXrrJKXmxVZti53McBCXEPTZk1hU52XeQjm9j1dhxKrrVMIsPZVV9
OmagF/jRS3rx8TV7Hjk++UzAw90wteERTqu0HqaPSdCj8lmskhZaRtEmEDiUJiiE
K/vIEPnv9lI6ckOw86EwtbXp+1AxTRzzJslixoewh6QJE5eO3ZVYm9It7QcpXNaK
1kcipoKZmFfpleywDwVf9w23aazmtvHT5rKA7JqyGZ8pwtnPYE2yTs7FxjpTqbax
IVolDDUopYzj/mBO2ah/Iff3S9buAYaCg0AV4rYw/HlIa8f5iaiMqUivZTT8MHLY
CpOpPEmoW7qgW0BaczGTODn+DdyAcCkfxeJfOBjaxmyQkErxMQ1bgx+oU0MISPvZ
BzS/e9YWxka8cUpJhKsel6rLR6613ZfST/c9k8gkWVc12sHP9xS/oGwqgNMWFWz6
Telg2sT9ybittLImrPBdnzMBqrKgypAYprQjAUpRoy38yxTO8PHAZ+3k6+CdxYN5
7o4Viyo5uNaRQO8SjvweXx/N0i3AuEhcbVpJDhK9eiTK6nXJZd0PgyklXs9e7HVF
NWMQiINkjGT/vj8vdR/M/BAWbdvAhzBGQuezDVKhB8zt9mf5jfmorFvL/f7bDXTq
9OvMSVUhNOgU2j6gXWlRDzzKqTDPWY8SVs0qFb6nold1FCNDzGN3tis3GV4aX/o2
AkWLNjUljGvWWTdTx5PzsqCbWhdsrrJZVuM1JMLZWwLgzy93xgL8VZEHsiYb2K11
3wfeb1JMEUXaGqqlCkQsaA3hgkj1UZzb8AmGhTgbLtdtIngYVSFEwmtud1QO/+5l
MWvDUMaqoHHcM2M7Veno0nLomo3WBPfE9F3ViHEnZcue7HQvcbmSk/rwc29h5cMm
8mMCCqee6fuXuJXSd7blXT5+ESJvTQhkyHp45QYI3X9+s9Mm1t7FdiHEbhu5DDJ/
AgM8Murfl0EJCsdSc8wRG1HV4Ps76IFBNeHZ55Ji0lQeRL6Bydg/KV/C143ZUQba
YDaCBdrIXY28DTNVApDL/EaAybeArQEbx3dyjlSPwPV3IboJCCGA29avc2aqDAny
ozYFLVaa3WRQlmcGV59BMzqCVEOf0sG4bH4Zac7itGgutXz3dMQR5KJjXBM+p1r3
hXq1Tqn4aTdAQbWyyFBmQU87XLU22Xt6pbDNnoCbikDUgV05QJlFBrgMYDHW9HWY
SfdqxMD2Vp5+ldmDFQgvzWsiuu5JVSx1eehcA3P001OJIG54sJQ45ZZkaj4ZeW4g
q6uGWdGF9y4Lgy1HaeLboPpJUXMyoFLJE9Vq7xhfhMiL7DrLSkQ68145HBM+evsn
poYKKUrEdYgLFCioz5PYuhioUJp0mruLsU9J7OMKiILoGlMN+/DduaiRTDrHMyx1
VJiyAlibld5lheukm8GtdZuMqx+PG3fAl8dUAK2EBZ96FI6GnwkVFQN1+pIBwvjX
yCqpzL0dc3kFJV0XP82aW4U09LR+GyRWb+xqrxDk3Bu/tL00KhB7Ir8BmUETzb4h
wsyH2gOIlZtYbEtbllb3sv5ZpESgn5tz5TnaJKHZCyfxoeHUEJFpqQHrXAQWyM7O
Nfs1sctDtZSaZlECTFQr7crnHSyb7ceRUtPpsZoXMbOieZYDmsY+GdNR/9LX5jye
283ixugtkIJTUU7ZP29MgFFth9BjbsJNmBLuAOFYgaMbdVI6tcZ99gIxe3VWITjc
hLMbadidO9kYU+yXNWMG2NzAgKM47qlt8+NYiG2PX+qgSX++QXrNX1RpOLyq0Yc7
xi0InbXOZ4zWX2Z6l4bJU4J9BI2dpLBajgMa3NZiGHlirDbnzvvV/k3GQG7NbGqL
IvVlJshYESj/9O8Xa7yHlmm/Hmb6a9p7E1Ndbmh22gWjJEly9BRn7ClrymkRugmg
zk7byeYgzM9+xin8QN39NEHl0gip4JrdspH6hzWIorqobErNS9nCLtvQD+AVbV1Q
1BBkWLyYEh6+2CsjVgpPr0wN31jpziHP8NqLa0832NwMIsGq4fqrOBQBrt2poxMF
9b0ooYLAYFa9M7JZzBXantiW7BX8QBApdLd98tCdYT8akeAQw/LYz/yETSPv4gW0
yMkQivcKTT6LSqkv1kfU4yeQO/6j+auyGTdpR6oN63MsnAFUR1klSMUqqK8uwfVs
H7A/t+TSSwMn12ykJO3Y4XsKtJoRaRIYiTwJWZdgsUmm2WJC8sl/Jsx5joET1eGc
cZpE+PR6CPQ+Kx8zRrXZU9feYOOK/F7pJGSlOOkgOdoTgSKb+BkzMDaOI7NU0evs
i/yduP8C7EL+EXQ5vqQLH+/rH79liTzX/t9XB54ndsD0/eHpMO4BWApTX+o8uqPc
sx+8ZU9nkoayak5lztABZKY5T9A0Fd2EGYM1U55GTfVSpVJZ9vH2s/xismvaEUpI
aJXOPifSx9G4wz02Q+wWbZQbLh2Jf1YWTkjyqc1aactaoCSKMvftBAjbf2I5zlOX
q6B7+i5FsQP6v1ZJppzcbCZdsYoEMeHDxFBoeAiCxD4sseit4eWWxpYKHMCLZZTh
TmGKkKHhb9gjhRCDVU12tv08BK+lef6Vh9bUOkyzCTPWNe6+M8vy/brrfnJJ8kc3
89Y/h1xMupb1lCEnY8WRPa6eriXD3RTKKTdzeATaDbBe4Cou6uUpZFV8+/sfwLmI
h9tQmlNc1jOViXy9gfNdvOr3OtqqSjtB+fKQZZ8RyPRl8AZwKJGmIeiwQund3LCg
UK7UFrJ1UK0jRMbXgpMge6i986HsEvI34t3SivwlWjg/0GRrTdyFauQHqFePDIE2
KbOJJymSYxCmVZyEWtydwq2ICuur4swq9Yp1g+M5Hgl+CPAtMmlGf7k1iHofRH1o
eghj7O6Uo8h1wVXPXgzOOJU5PJopIuwf2PtErEKlaN2xv7l5HglqvTWrdap1scdk
o3V+g8THrQEKmeqvckrpz1/Ar/vkwV5t+SVyK+iBMK6ExO3EO9MW544a/noyDr7u
eb5oN8LiWtfZFDcR0/u9YmTfoUMSizupWd83FPbNkyphMjxTxKYVdx1GDDy7xnFt
ZYZslrBciwjUm8ZN3AlHLQHXEXzta/fe7I8e5c483dJT4c4xNlINLKFkv4PQn/fo
1HRN9YUlDDcRe261mNTKdWwSCiJ/F5wLVotjSYsmLq2iN8pLUi82fIRV0ydnhOLZ
nvXGbtNsFEOLp6385BfrAINY2Lkef2AHW+NB+q2g72B5xvQCi08BV4qp6Ikh5718
QNaxXs9mxZzoOjETr7nevM52ouj+BD86VvmxP3lbf2vDoCBQzPmP1vaCj1Rs3ZcS
8cxi6vB4S3HYkERLdJoWpVbZ6QRV8yX9eUPfThBoZvcArfgHRM0OYy8T6TQ69GyL
8kk2TSAtOP5NmNFv0Hat4k77XdwSuUMJmr8JnTaR/Snhqqe071y2+pTFpZk1Y/vX
h2f3iqbN1znPczU8SSDUhcL/WV9f+7Uvtj0mT2OhyJVCnaclryveyZEPDBArTh9K
xCFwvu8P+7+sG7saf4RSv1ZmtPZqAiI+cCiv+mdSaLhSyFTlvZXdKdQ1/FGozg+d
PzInF0pclcGmpMSh6Wy+SL1kUhBBTcq5Lrvrlvec29twWqJ7a5TQUD4bKvSzKgem
97RXx3gse7ZalYrqZdDUHhv727H+jZbkXDOE2gcswrj4x+1RmiXqXr29mj2QA2tk
8B39ggaQ/EvpMgxTZXZTqsviK8wnJNxiZnQPMNVgFapypsScWcZZrr5b1AWXjge5
KHob+kbzLN5zIuvJWbPoKnh8OpzmAI8l8Wj7n5a1k2N0qO5XQkWC5HBCUZ4dw91o
z+ZdwUoptvXa/DjWC3NDpjlvQYcBAFW6Vf8thFvgdLHUMBTFdWcPLjaI9E+13u7q
zMQpgvbSo7AMpSijZ2aYT62+lanUAXa6TrJFgLNn3+AWj01awqCKubORvudy8dr/
K1Sb+zdByiSujxxHl+E1gd9sAOsPiKYDeXcKsN2NVFbBL2PxHm4rb0tipGKqPpxB
N1cDradz+y9GYAiJXqoquhF7yvhgUKbts+ieJ+WwAjsxx++ucu/mPnUgYmukpo3d
m9wNSndUrKziXludmlPHvfijWQB1hxcmAxYH7wN16wH5j77U6uoBZXwduk9zZC2k
pwmu5LLWs/UOAw3hniiEmDum9Yrf7phhdH+hLt8HmWLfQm3IK0lNfFgi8R1R5Rok
P8/gMBqNL05gUaqujYnpQ9vWaOuypYXujAH+bbHaWpvHOcf1LEP0Li52NANVu0K9
GFu8MixKqfW3Q275I+oqjxNixDoummZkIwHBOqJkOKWOkCfPqdGExBtVw9/DcOq7
sUOuiMsMETiPCV8iSuYqOkjTkzML4aN8K49W/9TbtTh8cjffF9bN3HnaPDsC+wZj
M13FbSR8IajIQcDb+JThny/0XDgG8HFjcw03GD5HOHCKTGBfTZYgAwoSULmmVcWE
+9LY6cZTda/Swgn39AsxF1df6pz6okQjqvdc3cnNKU7h9ZpMOaR7dm27jwz03Um/
ISIPHW2ly8yQXUfa+Z4zBUsmF1PQAEzdb4kk1ju+dOis1v4Fp4HydPbVaFm3Gcbc
+RYGjB5I6kYZVgJ3uWoYELejMtP/0ngG4RVNEphslFpcWmG1C5ysuF0jmopZwL4H
i65Yy8/WKK+KlUTdZuNnwQ74gXxGa27vEZM59PUBni5Gt4yhBzpN4TY5KiN0TBdG
8OuFcb0Ov3NpAt9aYFZMUfbaA8Azz8EWu1k7vx6OQNJOfsfdJnELwy/3TZIdCZfP
a1VmbyqrX/QNxC4C+d2x9mNEaNsnKUSKL6P9c7Namu8TSelGKc/RTbaaneDsmCVw
IV6DQG5IypCJUZCJhkFmlcSQAK2SK1ep6aw9mf0M8uk3+QIrbGyJyUIVStid7c2k
KPBj4euzQhuNmMXQCgcYKsmBEzeLdIIBsvC4hQFUquewRyxegxTMRPZINujUp86g
ID54PAY+OVaRmX+P+v/cQebz0aCEiWjzziSOq3it0rEVT8dXXu4Ui5b3Zmg0Pfna
qA9X20THSzZHcga9Iqixqtq8BnGnV6gVRKBcLK0njZ+byAQhjGADqQtGreREaLB/
VjPeHRBBqmM6DnSxdzCWO709xUMAwua/c87e+woB5sbKKxLS6mVbsttTjF1AYBVc
itWMhRoZ6V+GtdQQ92Vj+A2SysFhrlFPJmCIqMx0LXv0wBdsaNqZ3ktOTrLFPbLk
/zLmBRP53h9iy9mqsOip+y5LR3cmNvypptcUxlC6h16hB/BU8NaZANNuNdUVF/vB
N7pwZCmlCvvQ+8Uu0gvZu7DxqLaQdiWqVE9nYH8Bpdgl1fPcKa8lIgvVGpexeCd5
nR7BfGYdrLXWBVAYKhvvZMJrVX4YvnnUwWbGHlG9fYh1fDZW0r38NBs+lNxIDEqH
jrMBH9d9KhTAKxwvr0wAWxazC8Teovc+b0gyVTo8Zx9Vx1MZ58EPwxIyh1aLYjjF
UFgvElcwCthR4sG3oXpw+t6s0K/QlSHlowyINfTjxn8KWQbWMkXS9/qsAD5c7/Di
Xgi/NFP7s0ym0rl6eJfQ0Prw8gYDA2IjSN5JYw8lUZuNmy0/4KWw/LfgZ7uWfO/O
yVVS/CtMZbOTdtROkYuIHhXQGqrJrZ8K0Jcvej+khSRR012RrREDq/lyG/WZIjpP
KwqtN+xO8rIKpoutg/TnKx78ETz9kgh6G5rMGHWKwAkxTV8+nzHPmt4GGi2LiSX+
fvEXqmz7KEbJUZYbbyeigl6g8FrjCg6j52aMUiefVFJKbbnt8CI7ga7/R451bG2e
UtZtzmHm/Jji7RJDqF4IkmVjlZXMWwc5I40vLofSg4dL7LKHiLy/bMD6HoM4rqke
GTaiPu8j4QAKYaci5TtLygzIo1zCfNai6J6JPVC1rdKpvySbnF1tLx7ZSt2f0cep
C7G5AGbRXAd9DoxT2/7Nap7qQcpbxu69YcQryv86LOiPMJ3pP7XWEJ+xB0Ckdyz2
tY6J67rfSBXdOUjLEC+lDUN56tf1Tl5GtvkalFD6F0Cc7Tkm5Y2hX92g1lowPe80
HAylL576rzSQf6Y5IKY2S18zCAienvaMDDiDCFibb7X0WAewlhwuFSNMcMcviuqv
8UhJLkud1RobZ57Yt0bSeklLXWUUwZTzVH8vdjQsbMx+UeO/OMHt269cpd/X6M5O
dVakZnpXTC9fz0i9BolZ2DgMfAOjfcO7Mr5qoTxTG2U9IS3PDF3ftGHUaeBntIG9
ffjtD0ntbEfFyneI9kUtHq90N+5gumqGB3PoEbkO9LZzK6Hix9wQkvj2UrbbR0N1
2QgVTdEvIs4ggLP0Nm002t5Lw9yDRdbrthxumTyQEg4BvvpFriqZJNdH0GyJnctk
58g3lZ+yxo9wvyfBlQuVH50cCiBUJcxxBvLkPxfc09+GIeZP5SZ9L1aGjRa3qvno
T2ajbcOuEGMxWIRX194mA54g1XO2GCnJGTwgJ7YHcDjDo7BqnvhRm1UHkvcWxXYk
kX0u60zmn9kZVFmBv+mJQ84LxSa6qWMW4mSnC65St1PodwK8K07tbvKckAQIjNiw
egzuyFnycWhIaUPYWq6unf/bTPSIOqYD3aKg+yMN96FL/JCcSeBy8x/ChfpeBwdd
gK0lX5gqiDqS8cl0a7ZAlnbNatn+IoQwhWEhj3NIZjDQhN/ihG8hxo34Kp1iWy3p
p+jD+6OX7D85HZaHqj4EQEjez6jLBQip3V4vpKKdwII3evKhU077NUifG7zlpNVS
9hvU1b/R2fzyfV40xC+O8pzCTlxwNP49Q3rHQtDAg8BsvqZjC5Gj5bmYQohjo+OI
6mP/kur+bc1cTp3sdgcGh6JQJ0RzpWD2BiTf8wLp/9e3Yihrkq29edCUg8/Vt6Vc
iWjBorVIcKht6hzEoPcChqIDYn96Rqz9FnTZwZbkP7Aid8kXtVYKRo5raAIMGDsa
EcBlhqUPWhpv8l6OERhbdZyLLNTZzGaLd0mfBwI6qpzmm7nBiHBO3nS6r/uZAQNO
4b4GKCatdcotdyoldBn1I+t7yEw8b8JR+gsDX3/LeTTOo3BYT+qSutVmdybuaQ8Y
vJhT6UR/kgtMp9AEONnOgOweBepzl77GAfmmZXhhn5BKUd+4+6iZt/7hIIxixTvb
VeLX1UfmI373jx/u4ORXsdwwHbX2lFjURQwpO3/lAhFwGhz54RDyfZpcvRbUKjpB
wjzyA1dKFVR1ImcYvKXgZQHozBhkXU3Z9dHlnUEM7W5DYbvSEq2fqOy+haiozaPy
a79TNWeCq98wTCtUTn+MFwU6y43aEV7YRSG7OKZs1LnzMs8yXsfB9IJr3+PHylJu
v/yxKJ0RHGuLS8xnBhP63VFHLnko4Q4g1SqPzyEGsBCyFAnvnwmCTkgDoTY4+4I4
BCKUA5TJE1j+ibyuQmUbkWiaDmQptgDAByQ6lz8JY/0NDHh8e1k2PqoqwTMS5yaI
38fOK19F7vGEGW0VvFMxe1S30kVIBsVViWSQLDontI4bk99czQqW/zvRN5doFLsk
MSsOX+A8pB38b+yfQ6MgP8XsOTI3wdm/0bYGiSZuS9NlQRDj4Nlq+NjL7LjfuoP9
hViV1mHYL104wZ6oxM0VyGP2qzdVDgpTuPb1m8mvgH8250DflF0diBt4/FOVo9T6
O0U8dqsv3nw/zHLHABIU8Y1rcBNkOhgtMPn2lgCRLAi7aC0bBI8A5ZeF6e9/B1Lg
oAxdvCXkI8efmKTQdEM/pWgzXV1iga+R18sv0vhewxOLZF/B7VExTS7Ghx+Vr4+B
RR5tp+x3hMsK0H1hitcGOFJfd+JqKhNyzhrGlcQEScnuAf9S+IPgDGiv6PbhuoqR
4PN/2VAhHAuqJiFTRm1JAtOkqJE3pGq6vcLF9NO6lirIs1cJQfP8weeBS/sZXsmq
bn1KVTXdcQ2t+hXjI+z6EKNs5gnoQprwNBN7cthLeRK16VENZdGC4CXGDB+h0ChB
vUtfWuF2wR2OzuXPS5I9QVB3RlEO2tcLKGEbvMf6fw5b5zQV4aBCFVX0+BV4geR/
drTXSTQp78AGpLhkUrJb62CuhfxiC8lfYjO43ZfCNS8D5pV0C+CdVB2fz4nBTY2Y
Ha8DACnxJq4iNtb7T3xXK9TgCAD64bw91P65fRAD8ybCEqE1LiUccuueaW+BXZ9L
g9A9EkO9feIcionJ5SpB1hEfo1jSgwJcGI/JysMFmJQ/Nf9aK6SDnItXPQTyzs9J
t3fxAoAjqbEMc5QmSY3a9zV9W4Zl69zDIMUSDCqGZ9xcp48aGhYoVYw14ENYOvom
m2v6wZMBgnHOHxV9lWWUzrab8ft+mVw8ztWS7jyiAeeujQpAt6jgaGRH1bc0eTud
ZYfAy6HnBzgTho1MONuT6rDTgg9vshvj7d0/RlcJE30AEEjv2Dw9t+w4j2cObpoT
tZYbuuNmLCQuu0lnYTg++Z4W2J1LZbhC8qxrbtAwcJ6LlaQRB36qkTbb29TBE9KI
NwTdCZsTmVkJ9aYGMDhDJWRjpENO2EPfmjBj0fhzQcScpYu/l1VMSpstt6/mvwHh
BgqOWIDz0PwpHhlHUAfwuH8A2FSTYtHWN7R5OjSfnY9/31VhKS3EjA5EgL6hUUsW
45x1Ala4TlsdhZYvug+yQUXLnNU4TUbZ8NkoNN2fVTdFWCj+D6G23KpPlVIp97/p
Jo7d07CE28rZNtmSRhnCuVJgQDisZ/WkTUvGCmXQOmqOXGIoNYsOyoeibCrRqcfO
YiY/VwTf9WIehQtZAo4/NMYKAdEMJTZy6/Fd+MCTXeItEAvOIt9Qa/VbEC0Tnn8H
rMQ0Rn8+XeKc3dBvjMq61JrORxR4vZPMmubSajPQLFLhN/lyI5j/1U3uzyDrGXkx
N4tkdmooY8xO4NvlV0crHmPUQ7j3IDHcU3NtF7twLB2ux5yKlukwVkdN5MZvf8vQ
yqU+xcug8buEw3SvokBxNxSpdEjgfNnYmjaW8I+KhZaiK7V8Xccz0grK2cuLlP9+
iqEsDE5IAtMgN29y12WMAqUmJJ1SWi4gnSCjuK9l5eIA1scp7a7YKKsCmBIB2BVU
PbLo9lgOJilFNlw3/pcuIH16jjFUlaifBbmFsLe45hOUAQSxmSefS8GRD/G86QOK
ANRA19PKyhxjJPm/jM3hZbrXr9K5EyiPjqs3gNm2xSnzuJwBi1buMU1JftdbvvJx
aKItGjZs09mKcOcXYRhR+lJgmZ/bOjcDJG3dtHlTjBLI1ihFtXMcChB6d4clYciH
EIo/4liLEeEk3B7wmBI8J2UE0O+Amif66l5D7FDVrR7+Ad+xq6arN7rUn5RJ+VDR
cBe3/zTrOsMbfO9GOMZm33Xwo+wsWL8XKIx8GV02HbjZN5semyHb3s9Gurp0dVYg
hMzQ2k4XSVxCs/1pYMq7Ls2KDcZNtJSdF9rUrO3uq/YjUtO3f+WwGv4U3AmxiNa4
BotDDw9Z8GWOSRqSym7PmCSmdrzwPTVhKb8DYlGwW5Dleh3cnxjjIYUYPKl6Fyxt
I2m68eKo3nkjAYPGLI6CtQReG9fwSTgIazLhtBPzZTCMu+u3Zs+SkEDdj+kB09OG
MzhZscdDUsIm6wdasxaKlJJOiN+6Ekal+gRI2WyeYCaReEO5NE53P/VZ//8yRtjn
qtc3XoiFG5+rzwE+nIKsmoWtZZtd2IvrlDE+nctqaeJURgDHwqazUtio1Y745KhI
tRsYFt/aFeAjJ+zQ5ixT1OZ+wTRFU/8vGqgnEWp1NjJNVK0Uak3dcG5V12dsuSyQ
jRiCwa5qEabSh8QuHaLoYp6XWb8brgdZwO9fYyjFbVsxy6JDgMfn1kzCRaRO0QR1
QRi94ogD7Hr8cRZiUy6TyCiItcp5SMvEp4rR731DwT7r+UMWlg6xBVSg1/BPt45f
sDQhdhDI55atvCt9jUD2W3n04Hj2tUYH1UUVnMHXAWEyn6zHIc7xs01ymuPKXiNr
NS7eAP8SZhwojS3ZDNrFHvGtooNHSHDeKeqQbDr4YLmG3wZ5q5Gk24JWaRMdSIZ/
bI180ZUkBM9h5OBwaT5qPTyvbrdthKX0pqLSMd8/LbkE2g0nqFiLcZXun6omReU9
WXDvf38yda9s4BAH18VlGweojknH8QpItnpHx+uVsTQ5oDe+84XUiJQHwQZClEY/
UltDEagWcflbYSX43bV8ORlaL9REJ/09Z/Ft+V2CUYY2up+HWBP/iJqJSUBAg6XR
SRpizpKb4zIQZTvqBLxb3OG8ZRuJeZead16uAJpTTYud1d/6KBqi8kbYH1H3GOiZ
/DgmLk4G8ISLm36goTA2tDM+o9AD2UV7caHesDwAtAjB65LrPrIHmQ6MyWWo16Q5
9fiiPhzm5el8x8C2m0c5b6PF4fREIQfUsUYA5tUEjMWmAgi3LlMuKtOQGtAmMfze
xtS1WtyhC9EtUBLmElwzSdmlgui97gD1S19WzeTITbEazY75ZrCaoXNitTMkQAUR
RvI06laju5QNvaMFXacQwgF0ELtMfnb627jUDIdToxQZ6Dz0jzFXuDv0by8PaPHG
AdY8/AxzjCMVGCrU4eTEtGPKtSnpQds7/KJhJiPmncTa/1KdZhIrqxt6DrBfnuKT
l9K34jRUhrjp2ymp8Iar7MQXkhPzvsRO1Dt2SiHHEqZvJkV3sz8l/k+B+thIl0Qy
L/QmPiuaQI/XhgmsXY4YjR2S2h8Jj3ArXzEMdzVw+OOUX2kQfNDhjkcuBOvcmm/l
TTyTjXxcBn4XRKNt46cPLo1/4Ub55hqz52+UsnfdN/yYyVB7w8Kw9C6HztxYHFL4
XgKtgQ08QnsUTRgHpl9dzxd4Wz1VrW+8ROmcrIrcvtBe7gPhxx/4cEvSWNkp1KdP
tTxxt0uD/ATWZhaGBAPQmHLpy9Wrd3zxC707+Pd1G6GMIrdTCdH+2avLTHNnK97H
wC2klwMwvy8gRow9TOmlWyT0zN1w3ZGgwf/QNF2yAoVrDm4eOI2kaSvquuRNS6Fd
UwcF5hLFtEjnXIeN/n1v2t0guPMkGqWR/CHIAcNtT7tdEnPlqAyVAhRsJxZ7zzyt
ZwG74WWhJPNWwvC2smoAy+Ns+MRO415cL+GJG+bh5yfwk6ShoTwuILBS84HBeYBY
A+U3WmTI1kV1Ttz92NUHheFQLSn+k+KDg6kd+h42ZHTuqGNTr9RjtHzqBBr5CEqu
eqSdlHydPBjdGsxNfOHoeZ7XcnoTMCIC/i1Af1pF6wLBP5zg8W4NV8loceEWxNxR
JUdoHtM75pQ8QpR9Wy7b2I4aLUXqoz3JpbtiztcUaY5YjT6jh7BhOeqYVc0jUlrn
8J2KrPjlS25mVGKa2KMqL1hDDutf6qO8MzL6MhJ86V8RnGFv3WA9faqLS5r6NVWp
sogf6BlD64qUE/P/+Y26TZ++9WBrlSe1xSkJlvZNcbmwW/0cbQbubO1CfP91Ac/b
UViv2ziQvdve0sZbWe1yKDWfRCQz1IrgPCS0ezBEjpdKp0JTpfIDlgFYGEBpMYl9
72HA32onGgIwKZWHWz0wtabHEI1JiewLXKkAHjhTaBg2Ra6hmZ5YkdAreMNTQc4k
lk4S+e2BkEz7XmBT+uPDti6j1QTHlV/9s63PmfJZEJRTCUi/ajUhMJPh/0wt5Ddp
kiTR57+cyIxViCS7VxIG80NMhOpU2/KfHCRYdx50S1eQanljlOPV0D87igSWhvMq
54b/LFTLTCQKQT4LwlCOVB56K7UN5KYYZIprA2f69jRoEUP2Lm+I5zyx1R3+y1JX
I8730c/rWUpfyjqHh5usy1Iz5xLvxoV5r8YiL3j2ZZXH0OE+qHVgQ+avz7jRq1dG
Lo/MoM3zKvp6gtdC7QeSbTuN+XYk9fFMYHvzTp4kD+FBTedQ6jA1cR9bPP74foB+
OVf0nsAOuM5nJwaLTr2L2JSlvyCLXMuFKZuIn3rOtBZV5pP0UFaNptKj3vdXGp3Q
9LT8SQu1DtOEnnNHc6DpOHNGhOIiZNNwTk4U4pGZavG9ces/c8TOjPJmQ1uWmvgt
fqj24jBfeHsGbRgetyT4IbO3JN85p17mYj9fau24JHdh+1ZpKXiTSpWFKWvlCuoN
RbRJe/UASfvxmR1uhogS9NqqzCE3+3mC3wqUmVszwcdycEHF8hB9WPkR9VYodZ7/
WTaW+LI4BOxFKfVa8guztXGCcaz5tQa62WYlsQOOIYTej0/wSLU9A3uVCavJ4+xW
CRoM1dhnlbjJ4Kd2lCwFOduCJB0qzelHrwOYLkqpuY75FTr9wKJ+b5xBlsIGFrc8
Aej2BkflPWrana89W0a7MCaogAR1YZrJFK0YSBw3gEHIyjx6Unvpa7R1PbUYBulg
IQ0RRJE8OmC/pABb5qLGiUqMl97Em4NhvMWbQGrqkDxyQCoKNSLM6fmP0E9to6lQ
d2nJNNuqQ+pN0MUf/MF2c1N93Huo9u83Cs76rbH0XjIhRPPS0NQd3JDV+juEPK+8
O+0p2+1K2Edaz/UhsgzDAPHbx9/bC3K4ca8UgCpHMEm/0s4ICyDVVVrUDSpHxTlN
jinZona5wT1z5U6uUesXiL6MkVXFcXOX0HWPKmf5CR4oEsvZjJESWqS0wu651SZ9
fInpXwhSdUpyGSQqQkHd/jVrp5DDTRefkaYKK0L0NEQ6YzEHlNgfQOpwXGVhQ6u/
XaGyrB9QVwws9kUzXqMO8cKJo07Pl3ebMZGKQN6/zhhtAVRXvBvZKO8wWJAlmOBv
xAvv1MVM25HTKlGaBcPn1TewvRI0pQ7Puc38Vgn+PXKdvVXM9ql8WummnzFoSCZo
rISNxE9qDyozA3ga57T+P6ErdxDuK/S3/wbO5xGdcaIfqUXwQMKtONhB1n+uogWK
2MnMx//QN7TtO0Jx/oXjfwuA6HJ7cI8P4D37ytSC/3CP5POo4tW98Zimq+AFqW4I
XjeD1mV2FMTmtQebkaav4DS9FmjK0vxB8AZickxjEsrTYiUxl1ZR9v3v9vEFe5TY
QgtVrukXcM59irTfMyDZ3CXODmbQCo7nP2pXfIxDYJOVDzbvU/p7K/FIe4qTJa3i
uimnJ9hWaX45/eDChbfE8NFbvmLzhrnv+2er8sl0veHv4cRxXyzf2CSimwJ3JVQi
Q2l9+Q1LXYY38EjAB/rFNk0+T17u9SG+OgPmQlkXmNtDpObd4s1NAC7nQwBpJSgN
v0cvKacVMW5KQ8saiSqav1QoMDVCHo1dtADKBfmRg94PtbBkKIfylvPfZeXsHwIb
/1gRonMkeesQdW+Wznii+XxY8tw5wW4lfMQYPbR1uIGtmQL5hhHFjgtgw+vk8bt0
J4e5+QJsqyNEbEtrEmcHnIj6N9YiVhasEX9F4IjBkQuDZG3Q9zkJo1817Cn8WUAP
2SHyE9bCiqlrRm+muHylziRS2k4gWZkfhUGFWi4dDHIB9AJz/puCiwpMgHUeR6Vd
1i25WLLiwo+DP0Ba0DlpAWWo9lm+o1UXaka6SCYUesP8B65FXIo2dwWhxYj6wqjG
6yAV+SpLNKVz3UJKQXslEKczZe8s4V1tNzt44dodieh8UkB9N1FhPiGea6xY0PSn
d3LSAlBhmXxoOeCCrRB92WSLQXV7SmW702AGTsHLlucHnLdHrxP06gkHPYdXm58C
YaW46F9bCF/tFMtlT28otob47K+kN5+wy/uFw+piVlFqmEE4S1GdYbCCcpa1WD4h
po0aKTmDgBqoKVBxhZhAKBK0nXyzq8uji9fxTeOVcBWTvMH2OJaq4IoZ/2S0y58v
FneGurAQPrqbiLJsLNVWS9kYdWEvk4QNNteWSYiATO/gKszPY4VzkSa5grKNoY/M
wxYz3EjsnsoeVYhBvib5DrBnDNy+uMrRphftZClLW/YHvFlscU3VE7wFNW68F5uU
mUwTq/vhZXuM/gb7pq1YdsvYs8EelJQOh9/CysjtMK9kRxxUF57zRPqmq/Uybk4J
UP7XCWPStKea2hzIBLgsBRRuPbVdJWFFY1PmCctxt3D+Xg3UBPBxI8kSE8JBDXlH
5UEsyQM1XX0T1Ot9kqSkGCKOSm5S73RIWEcWiqvQF7nac7O1rdKNVOGVijQl1V4G
TPE/PrvpbllJ1WK437Bekgqx2DKq3zNloMuEG0wXsWxXZYVfJN2ekNz+XGVEB2fE
J69Qn4BHHbyDFcCoGZ8UpcY0pT7GmP7riDiFkAKHNHTcECf+Fz34DbCvYoAkvyEx
ENmSx72zMdZohNtUvCqFaDPRh3BmalR/GvUq6EJBwdx/WkGmEKB3krG9KuJJGF5J
h+h5w2gbrv/ETMmu0LQgPVsV+SSb35Mctf3xWEum01mktmOlIsHw4WBE/t3QLib4
ES48kUwRq45+TqXR0jCB37FAg3DVU+GKV0CiwrjqYRhUMElWhah/Ri8S4Q9WJDHW
87GVYWjpnnfnSI3l+kJ6Bw7pWuXNEck1fl8iPN0USsI16p3C/vCaXbZ7EoKyqIIp
x+4zCbQbaR4AhXjK6euy71iSI+uwdV2Se49p9k6FPssbKB078R093OThgeUjlVGt
MfLcJjYp53WJZF5xhvfO1SHatRd0IPs3JWCIfX3YUdwa4DVCV5R4LCR6mZ6v0b+B
hvfbuBTlPwd72DhzrJCsBr8ND1dRPotRV9RxJI2zEwzyLHRXW9IoTzh7QznCbzZE
W41269IP07OjO4CDSfNceyMR82MLfGXnqsHZeaGJINp4rxIYAZcyk6TUNXe6pzAQ
raRK/de/JZFISL/LlYuXsI6t9BFGpTNwvaD+SyEN7RVAzwWU0xOsM1SXNlnSUaOw
Qyu6cFoxZQnT/dSAkGaZLawY19KRhaiMKFA3IZZE/IRsNawSoE19XoKQousCi7AY
p4RvpzgQYt/DnPWXig4D5Ohqowtx+ZD2IzOlpLvcgsrkm5vMyzNT3NiEiwX0MYBK
ZaQ7i3R9BZ0K1XF+Ik7IkwJeIoYfsf7nQFIFUcINDihOxbKY06l583thdbr17Yz/
X8EwtGI5VWUJ5ygi2h9YfVDStn9qxGktHOLOS+8j/v3FkEUYr1hEuPWJkAbYbWee
x6j2d6U6NFx8u3OZtIAliufGmMXkm1C+TatKpS9Q5t4OAoq4OTXjtMoqHdUBiJn6
Kd+gEABG5XnBY1SWggCnBFHsYKvR+7f+Vvnx8ylBChUtqCqMlfAl5f6bT/ZVlqvL
jkMVBGunR63Z39x/ERimwcH7kEaVUY5/AJ3Ihf0UFrLBLRD1z/yBox2L67D5XlCn
YZ3XzqnsL2w/vuDzpzEBkGqqM5XWLL3tpCNYCyFFb44EeaGbxCx5TVpMD0j8Xs2v
c2J0NiTHtGmiR4/9A+d5v0BxF29QZMG80pdziA1Lpa666MEXd3ylwKcG6FsvtaZ0
1u5g32unMJVRs+EqFm3c4x3teVvqdOnmkrdrxJBjeGE8/fPeP4elYDvoMEYSvw7+
/INaHLIEsa1hApwxo4cxe/9cgcQnFzDvvq/WGlJkPIWOQY8Lu6+dx95+D1swjJpt
9zcqa/dm52r5qZIA7q2OYQ3Kql34RwNOwoleVzUgfM2vrOxw23dqrjyKcsLER9vL
1LBaYlSaZwon7b6r5vES3Uz6YbUTtN/Aal9J8VFWTAWJnqeggjrFP5E+UZb4BKoR
biHJEVI6Nh0VtZespOp1DpP317LtxiGhS+islwH4i8HitRGItEBsTwZJLGwO+PmG
XcHYq3msui5DP1HYqkegWc8P3qjRj3jGfFVGwfaFprsBo1eECLOLF2tEhM/kCzea
EtUOn+Au23qZ3IFcxX5EWIC/LcA10hjRleaT68gZwSrNUUYEHZxWBaiuSdid6jye
YVB6kc0sU/LopLTUxSOXbFBVcO2Kt3LhOqYCZLSfmLq1XLwVWmjw9YTAcYZ8g+e5
4dquy/6SRHgv7ysF198/k/v85Dqn2D+X7i6KbffoFk/B4PtCQeFimeLS/Zi1jsFQ
EsTyu+iKcaG082kCFuDeZX/jdF6wG+ShTWC9L3VVzEO+z/JbXrcwp/ODmBaKx4ri
IjV6U6NLNjgjkBMlucSYOb5ufUDYwc4V4HN1F1cc4z2N8RUUfY0xmzznkB+5rNGV
WuRSRMWsSplicKsV+wdQSHZq9JbTMjwXRK3ABNQ57xmnYhWhhqTo/uYv1IlwSnCa
qqCMa6OyuvsFLISH1KDhXMIWd5ErUWwUJU06IBH516HQI7j0p6WEPC6ADN/lpjX0
Lr1yprmWLMPaKX95yr7rhj4R8YcEZ3BRY/ysK821xYlBlw49Mk75m+jijbmWQprS
y/vWYVtCV949P7RysKB/gS/CQdk+op9fGkXyjVbpgIGS6+1SHiOkOzrndQSBLddo
ZWMnKUGss4EalBPnq469V94gUjLBay0UQuP5q1UQhmQNE7TAHB66hMghNcZneOLa
B8AH5wWOIB7orVH0hl7jO9vFw7E+/Dl99uPkg/TxGvZnsgNTUbFkKFUMCVYvcHl7
CAKbkLhVmgkJhbSnXIlbFAL4taeC0+CV0foJasts4PmZSGaEmCD9B3DYQPxzAlYf
A+4ddAZGac8fFFUhv8+L0b5ss7UHaEiLsTMvrUW6IYOFPcznabZR1bT6teZX2Nsd
3j2Zhm0ktYnFaj3F9QeUAOZp4TDIegTq+NHgA+2YDIBfz22WkKCy8XXGYNhOL6I/
nCDBtY6ir++wX97TDIdh004U6nCgJeR5xaplr1n/2eBcmTrxK+sExbM3X/drV04h
Ok58OF8xvrpKdm/k/hLtAwiHZGYsQPKP5IjidGOWVBA5LIR0gD2JFSf7DE/zBRWy
UZz2/pi/01PEG6DJ0BRFl7BSPEFKLuEh8VijttKd9bkOEgL6VAuc4i40DA8TJ8Cj
hV9mpf/yvaboS9bP6+VW7ze7bSJEe3tkpYEm9vC4zprf2+ZHweZdRplIjRrdpoZL
Zy2hqWW/MTXr+rdpXc2vy1nMB67q5aDvpbuwsK1kXfRhLriYNk1fhu96g01ppy6E
nhJTW+iF8kj6JacSXByCFDTzx3GjkHWOC98Vwr9r8cT9isBkUNAzGsEUGLzc6vUq
cYraj+1UM90asJId14hnvTpWTR07uC/PzKhiO35eMQPyyrM3AgvEgV6SCX1qZWZ0
3YlZdM88y1UBXp2fh1BPhkMQPHB5Rll8bO102QpHHAcnHyymsrMi67lT9Jwm/ux/
mJie+EZ4lu5HhwflhkBy+zCy3LJO1L3+duuBqvClqQ1Y/eWvY+nyQAUN5d7nYeUQ
nEockBljEMNujgPIj0Y0+oTldf1Ez7WoddvFm2bV2tm15YX/nBKaEw8U4Kw7WkJw
AkL4qGPcIkMn3u1EMVhU649c8qy9la7HUn6l0ajeziMtgTwDR3Ayw2nMC+hoMc7n
LYPdhI+MZ2vGO1aBc1WRLlEIScJQRC7e0uUn9QAbx4nB19iC0GvHHDw45QDpwCi/
f3xESWexU4CwsClKLZLrYvzLTrFwzVQwX85ZhM+g64rbNbcK6fw9B3JVJnGwKA+5
614uYZbyqVaVslGqG3iZ271KveY/1RPmTcA5C65Kp78Zp9+ASNJEHksKdft036Wa
JyQoU+ckJjpzo/uVHLh4yfpva07rK2G85lnnzXYGn04FYRRwSEGqr9RAvmKlNRns
3lszKGlZA3UeJRPBoCko+OAL46w/nTn9lmlgHMMNtrjEzE++fXUjUxpl0EUuo7Qc
7kwxGDJMdH1E0FNh/J4lsiyDr//5u/7/r1eQ2IOPCp7AW54aS9kvNAmCA0pfduvF
aq5NfJaesftEVuJblShh+ZlyoDD08hT/MP0++PQhC3g5pdRkz6KVm29Zs4Dii9QF
bi4ZsEw5k7CZNjmNEpdbBQbbOh8x0W7fU/QEyAIjtmG7OkN+AlAJKDRpEvXOr/BP
iLJXUpkZL3KmFngB9IYd+c2Pfmb49aKp6YDn6fMFTUVARr6vbS2F1SM0YHSu0vi+
+98LjXzFpZvz9BJGw3/P1eKhTWfNLnBSMXM03URY3N4UZPqo/ChBnN6pXY1CzqTS
1Mi8qF63DOQmmAl/nLFsqMG+mvEZsGSBbnglgxNJaExJ2NgSw12uEhSDULFBuDr4
f97O7ylNgg3w4KlD2uqGQGQTW24RvQez6bRA7iQAhbLIYtSM2nqEn+ZOj1BylgPk
UV0NApdAPJEbR9whOkYDOMt8xaH7VJZ+GBwoATd0/MEhamAUeNl7MGwc/WObWokW
OPICus+sTqbadr403Jw9Pfx4XiTqqAQTBcVHetGFz9LuUMBJNhVh8+aTmeVLGtHc
I8D1VtcddrfNCxNHNK3ugTLYMojTPaqTY1DYsuRUuOxE8ERBM4VQ/q8jY5YVAMR0
RrWWB5r1EFthXnMYFCftiLNAcEP5yEl8ecNIjdOvMhHipEAYkp5gFW6yj7eUQ8Yn
oPJlJwXVHTznnX/EfCzS+uBVRBZCcp444oEPW3jbiJueRxMC/aMwyibn7wV7wrIw
O3BNEyUtSScNoNA65hlvFedg369XmUe0xg09wtaWiJzhSVEud8YQAaFPhloQzqfm
ntz6+pvh/Mov816dR+0L9717uHQF0qPytpgfbe9wIu8lJtzc/DHKfukY4zuZ7QUx
Q8xcCURGROVBbcQD5Oslib1W6BHx6s4plMGVxxrnT08B5IaBOy9AAtcHkzfLT8D7
P0DyUEgKf9UQV6fkyNJ/y7Lq8wxPi288oKW/HtHbOXVzyRErfVeO4W786826lMU2
sHvyhmOY+SjTSD2BhnZl+8nps8s8oi3Z9wZRoO1msuZ6e0tjzubVo3DsLoFnJNDV
kvNJ9TeguhhLvj3FuyAln6Hd0oL2JEEOSJwbBMKQE0Z0MYkvet0fPqlzlBuJ7F2J
ZkY0fxZLcDnQbmrzNowol0pmzg7AfcNNf9VPXyMTOiaammXm1ID7EMyFhb5NUJ0Z
77bFdrEhIa082YNpSoYEWh96yHXcF/fe68h/JEj+ZxttuI7s/rNFx28xVqDTdjAz
Uu1LxJ9408HBwoEBakp7JJ3hKVUSB1lHOFBafu93dDZI5OeIcJ4xOzsUWYmWPLlW
QFWVn8iy2sfQZYSCUZ3XCXbOSMmLfPklx7Pz0j/doW6eG6c5R1UJQPSesyYluPS2
ygvMqXIALv8bDFh6pPboeYj2Hp6pmYAChmxVrWvC0tWwviuHS2JcljOwlk6pUwch
EHgsBYS5OL8xGn0lASh8ZMZIkXjNyht2qokhKoUwtdWSB4X426y3ADJlWvwgqwZv
M8zZSpuocXaBUPHMyN4PMrhoqjkxnWJjHAxiqjaPAyCRxCX8ppVv6CNa7Cpei3vG
x/2xgyR8s5sHQbRusyTfEz+tKHA46NgN4yF2Z94B0obpTlcRFObKWU+HrI3P3UZo
NvHu0rLrnNQ2J4Poijc+vK2bUkLkTju7TQS8SKv3j2prvY/igNtH+QPAXSWJPtgo
tX+E1ijWTYeJanarXWSiTf3hRZnbfvymqy/9e+yPpW9REj6boijYlcAh512T6TdP
pvP/uatXBJr6fkUqboWRCFeX43Hk5b9+DYd6yLY38B7LjIX4ZdCI02Ky3HwMG/pM
R8A4rVUHTBoOjp1ivBDtRkQB8e6TBeHMaFUfNO9qd45NmuQdu/P92XYTqeLVKtAM
hz5deldYbHXwyIfwfKb3wxkuhe1jKd6FamOPfc3LTGYwrsvpYRh+eVqhmGIK2Dl3
q3FTUqThtGd+hzg1nIx7+wefmAB9PJrhQ2eru3uyfi88DF0199LouPxqTJe3Dt4j
pdTm2+EPCiu+WKw53hF1HyQb655iiZCkaUu8lJzTDT2rWLnVXN6pKSDTlzCpWt4d
9FHNHBc0gbqo9cplcdk/LiAijG6f9YuPTlDj5zuUDNWGstUDm9ID0CxG77AVf99w
wKwhg2huFawZRa9rQ5E/i2ePDlOOd6A3IytS1gdrBw82S4PUp8OxEpENtEthRenx
XDNr0AZVGNtywa40idlPHLwZdbYpB6oZgjVyu+LTcteEfIFYJTDqqrtctrvsn2FZ
X/ZHa2tRDu84STiYhAPeilKi0xX/lMtCj+ZNY/32jq5tvV2BXejuMZD8Y6Zu6Ub7
P/2Nhwkin6v8n1PEs0Z8w25EGoIZOpVeTigALNrlWkBN0MMtCFBlt6VS3ntn2Ci/
fm/rI+E45rZlSOP+5n51dyQB5X9rqQFinJhMnleGoC8B3HVaPszuS1vxAyFQmLHg
TKtT9R6k9jT+Iw3fkG79lMGxrA9P5UlD++1DHR+Afbn4NQtjjHFdK5UFWwtZQbmQ
Wm2HGtFr4nbCTNkNd47HUXDYGKoXnByU4R/33zLFpIp5yxqVjY5IkdZzbikhLqzl
K0KaMsoqNFsMlEgilQ7rL9zy4wUGlEJoNd4pbpTdGMK7WIL28z+JlHKx1MU4QcZF
/oGJpSjGzq8nNo6npAsqMZZVAO/+cie3xYtHffcogdcIFATd9f5ulhgxhCJ7LvbX
q+e09g0H9kLc5UQD/b5GxM/Jw0L3/xwhwU7FeEkdpyrIExzxDcRh/jRQzrKZnOau
8jGl5xiop3iH+C99mFH19rimJLs8CmZzSG+w29FztImPFqLxRikyc+/kCqu5IDA/
yN24bVgSDPqPnGd21om3z38Ko1F18qmdpuwo0QVhoEfK8R9yIBPs9GAjckQ+6tpq
uE2SOtikx9qXzHejs+BcYEr4xhY2AIJF5xx6sMzsno9/8hbvDM3cDpvJPF2ysy3Z
XNuSK3bW2jbox0C9ny1bMwHVgHiC+zMC3R8uuckL7gRtPexz9Ela1IuENLGhPVGy
qDTkQrlCHjm+jb6BxYC5hVUhPvJvTPEny1F9jxMrrlgDf+6S6yld/vxlXRHNbSpI
RiqMUbw0QUx5zt7UhCD/zfm+OLUaHoWNzPcus0J8d14h7bXopXS8Ki9ZeiAEr8J9
+UYA77knst34PPrT+5Ok+//HqYlRerTKkKtFRTXmK4+fQngT2awLLenSrWKAaqRC
m6P+PGAa9fuFilXOTDXs5ar5kblctupm33pKvabeXAJJEmwEQwT89KXtlq3LMiR5
jMHdXqp/4VlFxE9hahFNeGCU52NSdiLYuOiFfAOBXDE5H6x7UZET1TUx8ppC/Gik
MeiNXAJYIwPCkaWBv3WJOcRJPpBPaJQPNqhijaQv3gyVIzd3UsKouX3qZhfqQJGN
6fWGGi3wFdYZ+xhTTPeqHxsnUwi7bssy89FR+6hQmnSH6ucJShso1qzORb9FAn2F
fiEO6UQhLLqqeVpXC0ml0qZCVw19s757T8b69+xepJ3np17AxcH+vssNHEuGPnWh
YAwkW+ag+OoqEaulEMODNezxSREsmD7laL2PaJsNqxIUqqgdFnrVZM/90xdFL8ie
3TgvgZLR+4r7SWZYheI6p3ZRo1x7UWf5D+c6VbAfnt7UMo7Z/R6EA3hPLPk7qdbo
mlXIPbQ3+yJmrJJwCluJQabN0GKnK1Vni32XrdqeyJyd5USQgmYTRX1VUH4ReBQi
zHd1vNMA2uel5ezW62AlZwbGe+37chl7NnVq/WzuUHyn/4WvjhCa4iLyHwB9EA9P
+1ew9mcgzWfhrhFisFosOmSyIX2o/pRjqqlLUWO8eZfzL2sdQ4RCcOFadLG40OqA
pO+ob/KJ9q4e7XvJEYDhm9m3iNZ2PFkHr2eHOJBpG0YZ92FPopFnFO+QWcSGw0FC
8crB8P8DtkfKukXeliFmrsOQqOl5/73c+8MhBanMdZcD9/Rj1Jjdj9ZG6nIj4XXa
63v7OK5Bz1lpLniVYrORrIzrdoVTNWlzqGcA2RKIgsZTFROA/Yzfw/gAtM6Xp4+r
VYGHmHewWmoQ/z7L/CIbgjB7jyBw0q+qmwWe5C1Ts83hp/jckSM8yfpa9ZoE6Jq7
pr05BoB+6i6q9CPCUgL0hcQJKMshb329GUT4cI11xLRlUa+IgOuSGUyPh7qUFyp1
gI4RXF3WbqrLF62qFqYKUTr76eHiLX8navsxQpHJFS0wco8i6nzmIiKst58U+/cg
rbhVw4MoSemOcEYb/wJW04cUmoaUJGWlYyLt9+gDNmkSbnAfSbhuLYzZKXMgA3Vn
bBqkieCENtnB0zJ4yL3IYwFBoRjdbyehyonXP27VcdYlqBRd/kQaswFw8XDNqUxO
+nr+YyIagCPb7958CD26VPfSjWCidS1ejwNKmf0pMbEwSH2Ab2NueHGgxbQAYQE2
NSqLJUGXl4YxeHlXjGjV5ATEeh3Uo5IGqyblCnmfhvubKgM2xoUd4q6N97FBiV1n
cU0+nxrN5g25w5z4bySGdpD4QIQNL/VfvtdeE/WLA4NqRYNZpBpTcDJ5rwJ45pCN
cvKipnfksCduYbMxritevIgZA0PsttP8QR6MMi5AJ3VQIOnwszwTm5IR8EY/xZWA
/qCpTurhJtDRRwCdmRs7n/wBF7YkPhLS5blDgLuVKqXX4WMWN8U7VTKoqT9geXL7
A7IDOWHjcP5cyWb6FLUMTKBEE+omaJpS2kKdG3Y2+NT0udztRwRUFIiS/FCUKHo1
Thi/rFNMyH6/G+wnXtamZiM7BmXjuwgGV0R0VVTuBus+4tqmLJFFByAec7jgknf3
EhC1Q4LeDHwus9epzXXw6m5ZpsrFdib+HaAkQTDq536dOXldJLeYGhcmGPGTs6Yy
g9OWcAROPYW334/yguGB8iPf87icJHIjq74/EdeUu3n6JDuNfjo+bwX2OWxUUeDZ
vKqv8f9G6dSWiJXax1uwMnqc7mRn2pHx9MQOg0KTda7qrcawB5n/uLJQFwDDp+Dj
iRqNt8g7Xu3Nfyi0dPb+7PzBupKYjEKygsWg4OLDqFVMtZj4lDOeYNtGkkVHGZNb
NAFpMI4wqSu9NL6N0afwmLac7KbEHLdCo6eHxFNHu6nI2rOPXD/qm06Xj5cRYtW8
D4KkYg3+Ga+FQxzmKbhU/5/IAcnp0Lf9TPTBUkfDfZZUG/L1sjLT3jgqtoTUcD7Y
ai6UF1tLP4vphfJRALrpqCtGzufemRBB3ExSpbOA6A96r2d0oX1ll5Y1xodX6Sxs
QX1thsQfHsPSVTZSr2+Qz4nM6nAdqT4tVq3daqkGbIpjzUE1gSr2xLzy95z+W2u9
jFFfrKIAuzOCPVZcg4Q/CPbkgUd5UCDfdNfLIFtPs0qotLuZ/5CgBDakNTP+H716
SKpdWr/0A+0NGvr1dPpiKp3o/3hcyEpxAQdT3DSW+CEDXszxVvh5d8IC5+3KKfjW
ljLPQR2JCUHtyl+pd20P0SBCMaEB2NFGw0WY89BkwupJWSo91g0a5yI720Q1JSxg
BhLZKjc3ash4wNcIfjbENLtyESJpP67raFdMWMz1JUH5OJFuPrEss0q8iifpEbOh
oc5grisX5Fis5peY2tQDzv3xlL9v/A3+2HnvTfhIlsLYiQWV1UoQsEKQjs+m2t4r
6lA+toPz5JGz8XjkRL+l3ciUw+2DqQqobjN6iLYuLj0m9IyATLnqQZzhP9QhgvDK
06HST4nod0CqXpjeAMYzPKRKFdB5a6NrBfE3XsDWtSjftJ7yBoWG1DJbLzmy9OlG
iHDnFbemoJ9M4NCT6wyAGLcDyWpz86F+61V7WtQm/jLGUv4y7vSztI/gpk/gOyZR
Iwpg4YR58Ahatb45fACJCI43n1TH11M4lhIzKeZtXEdrvMnC9fmpuy0E5J99Z4/t
pCB1kMS+Giv3JZoEuv+WK4E+7+fqq7M8F2nhUwnRiO5RMFIsZSEiiy57JlK9wE1C
9N+Y6mcJVJG3w/Da+/4H7eO1r3fCj7jyZo7JJiWV5GFHKx/yX79q8NaQSaIFg8fK
LQUZDqo56b5wdkUzWPSUpYFEAsQV+XzQIVb5NGPZA85HDf/HZf+s539WglP5Pkvt
HiAuzrnmzM4jmj06wCMx2ufip8BgHyCCbm/4yMeSSJfMDn/eBe9vUHrMD0AWSNDp
p+JZSvH/CsiKWvLvJFGCqwzKBLjKS2qcevlUN4jhPbU+wGGpfx5/hFYykUaiU7ge
KIQgCy8mf5/GvL08jTFXBmL9kwjqVrz6LFesf/C5OFExWWwgslz0r+zqo56AJtn/
nJ2GP+D+Gq1KQQYyCcaMErXy/VQklCh2YFuXOFFm0JjqVCXD9FSmrjPeUFzLl4BY
cBFXXRkDiMymxa8LSFZkZSS9GOL5DPUWpy0seMrWHnNGGxLAMukpiHKFrkU7lf2D
6bsAGfWEfoGCH1yKltBbgU4gE8wN6kbi+Iri/FxGThMNMN31ZNdjIpYMTNLWzD+E
pqzSSpFylH9xR86EkWF4glUxSU4EmQUAQwnvINgd1Kj3JUDWqK/JylAWEEUu+8JR
/S1nki6DnnT16JKoM4RXMG+DAXm8qnRLntz6wgC19y/JifHshih2Y1iPVnSAB+eN
274++s04JivkFkhAKS45AO4maUaYNBEb1ZQRHjyY/Rg1zYgEb4z4QJEmIHpZOAg7
tJDZRtsGZSvwNebg4BuuVqIO3PGZASb2ELc2/R9Ks5+9hdwTW36hLCwjCkFEPARi
GrKAPAt5/GowLrpafn+LzaQmJw+8GwM2Jzgx7am/UZniwok8EGbOo+Lmk+QknNbV
BKTDt+pVaE4an1+GF4ynzgKqpdzPZl8HQ9+sgTDXHgOL7ZaGxBzY5as3gzLiDLqo
Pn+lpIMXiFz6Szc+tXdf4zpp4JlBx5Q4eHEn3NqMWpqqkUcnWCOA+Sw+HR/aiWEm
W00mNQLxwJEtK43bBdbkBSMnEo19dyMQeSYWFhYl6oIz/m7TqggES6lUHytGUXZy
UvF98sGK8JCOWIhZNRKLgucgtPBT/cGxwZprR9UhUqVKtE7lVfu9cAOEpCB/wcTH
tfk26UjSrx3ZNNdEkXFslJ9esKvWMfLvCM/FudIE+4VyobohHc72JDKEw4HkrV7q
Lclswm1cyCMe3D1vywGmZO6tKZR/X+Yfx+MfJQEowyMwcDahemFYGkM0McdRvy31
mZ7l7koOUWP4oiK0gMBxMSCGGEpvj99rfonoQEv5ASH4PkDuG7tqPUJLO+pIAytA
SFck7ITzgKApjQBLyF+p1HTe9faUEfIz/bwQSIihAsDaJ00eEoNNkVAsArLAhCy4
12edQ/8O7WOLp0m5IZTFFkNXVdCzZP8xpC8n+OaFGY+gJxvem73GovwsmJjb8+lL
JhVDAlcrBuB77W+g4aWu9aDA87TfyQvsVsiO2N/CCGSw++sMLLO33xKfo6ZZnOTG
UJ7O7m5HC1WCnfI/BD7DGJtDKLLuIgylXLubr47oDUqujryr9LWdfJ3QbyovRnjr
7tTJ5W7J1daAosjmiU4C88bQ5TjMFKuoZ1AYkBX0rIO9kYlym4uMSJzweqMwd+9M
PfczjYAm27Urm9nTr3T8gJ1yg1RDIlXjVdfUVieGeiaRgLzCWfNqz+AQwgSqFn2S
tjr8AHjxPiWWscyQCUI/brIJMPP4kqe7MkqW95w1ySVZ6U51BQnicD5bNvYvcrKF
qxu3X4A+k6972B88UTiPSEhuTTVgbqy7qD5BpgIoDfA2T1GCegUa8iZK7wrjKU9F
XdB01hgc+HkwaSXIdMB7ql6hb3SE+nh+8zbF8nQyZZ2QPYbaBIVOaECoa1hupto7
8HpSNHxLa9Lsw7moNzdIMnuZzqEn4NdrxVkJv9qlfKbz153iuO8ck8rCyVSIkifa
N/T/afMhL6/nr7HYg9xWNCh5EGHFBSjmBDsK6TBkGhxZhjmSQjd9+qPl1ZrGGBGz
AiDPWS01nHMLynRFzFfk/26Or3nM6AXEY9H3o60NW56HdT7+8hMI3kbmnoNS7HEV
kKpRsiHMJREo/UuWiLCqLGf6InBpX/tpEesyL6kQ/PxW7f5lnxDe98waZOvtcv7Z
58UF0BX1KPZzyPpptNd+yFej0B1rS1vj0bvcNXFScwVdUDesd3ikRqFazzvcV4dJ
eCHv7LAZ+LxMkVclQjhexF5rENezq6w24dpl0x61cv5qjAphiZddprvz4c58Ity4
0kfFCtInc31rBVJtm1Qcq3wVlw70B/FluTHI/NSi8LTzHv5zvHs25xM3NeNro4Kv
D/lMWo9LWtjQQsvmDBTzxRyWdvEkyfCHyMaWNn7Y/pnQ+xWsPAVA0VLE0zAtl/H3
1+4w9Wam6b4k1aBJS8vYhZitQq2CXHvnwxsC5l8IqTE5/rxC1bJFqI8u2NcmdXk6
FrrxXxYQ2cyV8ElMNEh9BXBIkEXvBT6CdVSe5tDCBTfdXc7yhBsVZTYlbGDqATVI
hQlOjxDh9PslkngmyWtAcaCq/o/tbxmrwWUxnEnRCulLODA018fztloc/7GDz+fK
rCxdBex8auQZVc7jzdLw4wGOO3roLYtTo6VJ66uTu2QGEMYZ+mnX+wBuDysIhnB3
K0sLp3LyZnvbPymYbvbj7eXjn5iKqEPZaurDzSsyUhAJsnGpu1nyMmmoRy+M8BFN
8Pej9ubXS+awqxEzcg9xWfwx79HQ/zAHQmYI67rI9y0KdqmMlPsBZH/LvQQo5PUO
M9NsVZxExFuhrLU4nFnlrhcp5zGpviKApmXjPQTivoRWCoWatDUEYAnSPOyOE86l
HhN5S2eO+NFI95FS8vr3A/KFspL0g2bDXAQh37MWtAX4dTCNOr/CUyhluQwgRwj4
/FcJw51FygXnFtZBWtMK74kw94DSVc4Xab0JR1LiUitSF+TSm7W6FECII6MslMHU
Ayryu+6gc3LXSyu8VO9TfimD4i6x0BALI6ir2LM+F94HYj5SqlxjwWl2kTArp/+F
+EnW9PU9jYgYbJ3kjntS5hNOUcqqDMyCBTzsdhS7KwFa2MZW2CaLVU6WquwBk9GR
J8MdhbQXHKre2PkqOmc1epwJf0nQJAxCv4mR6i0rCxbE0KAhKSiJ/fZoj52Ir5H3
HnTb+DR/kzbc3TN4MCSTEs/eWt2K0LkQfsaqI46HA8cGywbvGLPHUR5WuPARDUDx
OgrhSYuXldbhsQgFylAQ1fSecJPw/14lXVio0YSctjifScSSCAIRAz12d8J2DBCL
1xe/mBpouEQn9Z+fjwzN73KlfUlhxGephG6gw0lKK9yCZu74W0nqWLkfD5muGeZc
Rxg2RcSLqHxm5DDpO6j+qnpcpRW1C+KbtDOfvzRkEAOuZBnRphkY/DvLgkLa9loQ
iR+c+4pqq6E7mmn1iL0RjEt/Z3O3g6Jw1LDMyW8uOohVPSULBvaxb1Q5fi6CwuTE
Vy6cqba4hfeJCfKf1xNAY5S9Ssx+2e32JsnOKTNUCwaVgCwMtmKmyGcN0lJNGJVL
DqOCJrclqgtbbvU/sqUSEAVwkzEpxL7Bj3ZjSZcneaoTLGJEO8ESzU21iWdIuPv8
eRxGW6aGTOvv3GTiaIg3nI/4chUolszMtfMASpI6PCQlVdB0HkpSyHsU/hty2Z9B
lAUNRFbnLnoVVHTz5Yo3qDv8Ry1M9BS2rc37055tCe05+QqOrxN4L2DlQXgUK+jq
7JelEKhaoI5YpVlmKK0Mgh4WN3CrFvmjQW2s4nIRRJAgQjOVfyeN1txAluCCQZla
GGA97hIb0dGYZYQRMAsYl6SrhD96YjlhzoUx+3kcZwerY08M2Io9G3Hi42JyNbhY
c9xqfX+F3TROmOyEb5xBnt0cGQxKXBj010AOyQPjv5eXgvbYf+z/Wa+7EK6CZaGw
iAE8033XBBf4DmQq+Oyb9pvj2F+ZhT9IPGb1xYkttCRYk6yL38kLYMyd3mtqyrT3
fm/p6UUCjLTlPNw4fK0cVaAFnYnxPBoNEbWxw6R9HgPQlCO71pNTgeMsZGZ803R0
rQ3QSXdX6xaXqgfxjPXobhFG0Zhl0KTAU5Ykpnla5AeTITJ49MbJhwtil+HtRVhA
79TQx1tOTRJB/Wa2mC7qfjEUnAxYjjiRgfxjU/aWcz5xC2p57Tv2URyElqo4qp8M
Ik2qSDaWPe8CpsQ/Q1/khU8k4KPo0OOMzuQaU3GSAmrN0Y050oQctVAFStn4BZL0
n5AYQAoPZot/Dc0HerUaloGa9ieziUajlwG3jhWWee+yX3DhxfJ1M3GFB1S7XzaG
U4+Sc0nxm5q7GEE81jyWxKC+ZkzPlbMalKFvDAQlKNjQgNfmDeOFHNBYh2B9sv6t
T2CI1iIoHOuIoyjr75lf/XeneHJZAwXz+JYdwW20hByLlJEfRMiXW7RM7U3Kqcjp
nZgbLV1H+DGmerxUTDNoNjM3EO+OX6SKXVkGwmxsGSZmzaO7Go+ZP2G7+2pX5zW9
R2bIQXq4cPl81WI2xpxNxPZKhM2y2cOj3n5gsnZ6PS/C0U5Yicju+jsNlRNOtF2f
7fksGFi3YEBOBhvVIP0lW5VkeZ3xfEd2h8AC4PajGtIz1FvypOHoYbETYPtJDTi4
Kw6yUQj3tWblVD6/ZhorGdPyV4lCTyMS1etBOgDaOtPds3vPOS5WnGxXhTwyAYKT
Ov1rd5NR2yDDK6h69S+BytbSVbTqgSNkDHt/ZjUQQvjNIJ0IqKtM5IQxRIaGCHjZ
leiYbh/mmTCVZ928EzEM5b9A8E5/0mFBFh5Uv2iOeego/bHmfh/5Negff/6Gris3
uTTTkzvfAvvfkszaw1UB8UErr85nEoITk/wnCsYAFDJwjkGXruV5+oHTglUKdpmk
rt9FXgtkU4wUu/TOuzfiFwKvMQxriWEyqU/pSdIf6MfCWYNSQ/xJG+Pl3ULxcd1q
Of1YGwNHe9cHPA7vXBpYODsvngMh+g/l1g0ozPdRBOZOhf8n3jw1obTN13gTja2h
Ar/Ypk+4PZm+ipcrmnPs6hzrZ5jN3aLS8/sC9QPMxWnxd8OuwSfr14KehQdWlvvi
otp7E32tgp2ZC56gSyujgZz9nW0++ZlggyE/KipZeSfaXxAXc5C8DGaMgrpolXrN
OXsqMbEG5LNjlxnD2dr2XWhjrrJ8q+08qpja8qgrKo7CQLqw24tokYYHYUUAb3iC
rSp7oYaXo5WsL3Jr+1o9cBw9hC7Z5wYE1PUH5qFE5ETlad8Tm7NxTwp2ixqAWOTe
yjrzkWmXk+1sbFKQtn2ViFlxgNsGY20+a8qyM2SPScjaV4bT38tjpacrD/3mBwdM
L7q4bHlRggM1gT+eYmn+0g818xdyYChretmfsYErDH5lV22TK1I9qo4/cu5BTWAP
ULNTnZiUHrDesUgb5lVjDeuD+/jFJRO/+eFaEzNXwmtfAPHF3tV0gTVUtq/SsY5H
UUJjDyGhL2Ba/VP8LwMrW2knM9EdPCs2r1JPJVfEZX+D2u++qstgEqFHgffHC4kR
R9ndpaNXkmppJ78YBh7+cScTFBS2uq3Jj+ie6zvgMwY4uDBT5Ux0TbNLGDjH7Cef
+5PcIrB2UEcFf7uupPn8KxbcbLExwXf5/BBmstjKwi8HvudwYu8S0WWntynh1joc
bT9RnyeB3plcZrd3Alw5EcM549mCj+0+uJ4YgVMPj7xhP7AHaQtTcz+fUx53cBjQ
9SfOqOlRW9GKoRDMXEZ9ZIAqtPtrM8u59Pzr7qTmK51Nrojx+sIb0J6Jzb6RI0Aw
DXuMo/9b/S84oN9nBVfFq41I5y97VyM0/8w8ld/iuZbU881LHHzTPJVEzYsFm4AZ
wUDB9WkzqkUwh4evo11KD81XYHATFjvTj8UTeAxrllNSqF2g2dF+QQNKyabvOjl5
/Br1/IaEjTSKPoFGcZFhHW1jrAxAS7Ku7tkpf7WkQenXKPIUOs1pqBezDS9jnlEt
4GfwJVwiIW6/sVQtgBR18klnl+70P4RfwXb1RLgkkciTCjyrn5AY1U8VfYmDziTc
nGMdF1zfqadZ6hThSRxbv+WOd22zzHEgexlXKwTqmEqK5etT8F1SIS5XFQoBnlmX
kG0kT/sF0opD+Ecne8anBHCkk4ZXFv8IpiS4KhgfJTaAYV/Ir6VoPjL0/kuF9zQj
727xJRt66k9YzAw+3Fxk8TUP0HDqrSBOLOBMHbHQcAXPG7Y/3Z6GhEJhibho5Z1v
mOI/cx04/gKYo6Ul6gCNX/0NESGKgc6628rI35m4vSSWBoC5BxToRfjqsHHNBey4
hzkqto+9OhknQw3PZUZP277lDGGTueyewd5p0vMRBN3ampDnDg078BrXYI9MRg8b
HqGyZkw92kOKrBRbaaDv1DOrOK0DUzyZiWR05OJ/HNz8mNlVzhX1sio8cuWoC3fA
qkj7XxM4oVIfsd+YPUOCwDeHeYf9B35wjc0yQLVoaoJ9DKce0bTjOkikJREmdeC/
MBKNv0cwxeJENVmr8Xr+5TSruPzD7tW1rtXPifKAIe87wOMv9pAJXnYuFmSpk0Iv
tO70wjpczNCRMAQ7F8FQTGAlkI5X723kh06BCd5Z9TeIFJvm2Jt64doGb/IzyreV
ZPkOXVXVSLcIhui4WQfcRse7cN5Dh/N8ozTtJ5Cn5ROEAP9vW6m8PxZ/tXtzvlgZ
isYXpyN/eSoaiJ91G628UiIoyFfaNWC1XEFvUp2k0Van5gaR6PZxzsYPRf0vchL+
GfS6+xmjoJwwsmG7DwAqEKhPGxNRQWLGnQmhalxUz3tsOuNi+uITMTN2yL8CjXbM
/m06a96Ml09h+S5d9uNrM3wj7oWZ+yIcUZcZ9MGgbJiGesD+GDMXpnjcsEPrCNVf
ozPAXZqI1tsm1OfZ4eGD8kywppo4IUv8xFx+7+YLnJTCnPJFBNyZXT8Noa6oHslW
m0SYDq6PKI9b4E7FAbHAOBfIL2tBCIQN5PAe4JFQoVOfgOxnKamOUAnQMiYq2n7r
6x2+pKXD1EMMYsyQucXFIDWuUeW4c8UWnOOqVlHpzjR08/+H7siMeNoH0oXJ++n4
CvXAmrZ+bmCJxsEma8EEX5Erl01S6O/6ymFLZ8WWbvVLLmxv08S2PieFx/yYhQF4
CW4pdn5kc+8XGij/OnX+M6reDBct3AiBgFP3PbNpgSRwxVTvY/DGYy2shF4D3+W4
kp97NicVk47RhmFY+WFpiARi3qu7VZiWkmCrGiBiJO0dITV9P7dmhd7ffYqWn4XR
sudcQM5WRjHyfS/SrF6tLkMTyKig0fyEDEk7aiE2gJIUIRdSxSi2GO7sNDjA/F9P
XRDT3z5Hhdupq10MKFl06IQPNncLJ4QDuYFRBu/V9wxm1tmE8eAweumwH9riwZ5v
ILW+WOw6RKp8u60959gawbA8WkSKsUpEKH4kHo0NAk1+sOPISwGwNAhsE2wWIb6T
VAR4RTz3wvCPekGoqzgcvspjhA9Zbfs/1HDpmrnOI8BDXoXYv/DRXsNRvw7tNcFn
o0pyBizcf0FoHHaAdIAjTQ199yoYd0WyEr6Qe8UM3PrkqymJB8V77DJgq7xfCIhU
mL3lB9mWFjpIPQjJ+613cB1RtW3bUFGEOHUaaVlh3223bGa0PfD9xP9ylsMhJEng
7ztCJ1kn+ZkhXZ3lCXF81JRSxzkVVLx+wGjstvzeKDa9D28dI/w7wzrJ9avyRuin
HOUvox5dn5+aNoqaE1bkDViwcCpjuX/oVpxNjKuo6NmNsNZuij+sVEEe3e2vzmVB
73femg2gqY+xiETvvz/y1z9uSfDgJQquVqVJD0MN4KSzpGS5MqT938fkzBa215Ql
K6Xx/h59qsqn/dwx91TA/jSCF11uA2ZJbaM1cwSgeWDcARy9/6g+LrdhPEuVOgmW
HRtu8YyAbaXrZJDO4/fTN9nvdTYxy8ZpJWZjuzZEPDmwpeLqFG2RrVJ5I8so6u88
m6P0OlYBI9QNVIyoAPfrvMTOeGGtXxGpPnro2JsX0YW6Cbunqf/sFIHva3ZWH2M9
EjgvT7F2TbsH06/zGnr4isS+7Ct8PybC75W4e0aQCVBCGkBEs8YB7YM6AtD7+ECH
njBVXiXSf2VNApqOQGGvwKpFo3eijjh199oIiIBVAy0t2CRREobcSPkh6yC/prnd
wfbYgInLdlIRu4TmZ5FFaRq83BZtl9thWs/edVErStN/HOIuc7ocrFZqU4uonynp
osvJBvW0gYlRUCYwfCrMx/PPlpfg2C0Pq0pgu/f86VmFNtvqJvzfHJjJeX2HLZsz
/s/9AJLIuY/Wa3IYsmBcyNyPjmRpfLJXlIzwjpPJ2xElGLisqMDkUoVLtZvW1D4r
8XCt0cRLaDhc/adOidtalaPPk38EANbD99iQozbPd+/hm0ehHjozUJkn+qGc1Fyq
9wPTEYnDx2Iv3F58stDbhBPCYOe/oWGayIF9SEvOqs4TlyrIMO3IP0PqjzN9mWJq
QZkN4T3QJCoYdm5dMI43jNoNr1msCBwth8AybndhmncHaVz11HLMov3tj5CMBEl8
O/OvGl8z758OrEhFJgfAQiHD2gISHEZ3UVByUySb6/GH4xLzpG81MfDr/Cvht9WD
/HQh9fqoi7tkn703x99eH3oFPBZYMUnU4rZ94o7VUdTNS+oq8lxooKVfWYk4uqXJ
f9ZLEVO7s9WQUJmvyWTNyQ58ZPCIplQUToM7Im+S09FS27hvDjfl2Klq3Y9A12sj
OgmC/PSC74WSohn/alGMVa0GXcZl6xIILLCzDfBB/jeQOI/NxGD2OwhhMb/Vk0Lp
BOUA9q1MPgBOpWqDKuahTP4rF/qZGXlGKAP1f/j8RM0bwK+i+UFP8+Ru9G3YBV0z
3jn3Ex7G0HaqyWay/My29fBVdOtLN/CDor4CLBTed02wvAC3StrsbwK88razOLol
rxdjYaYgAjRxgQtQQ+05X3v71NBDcAhLR9tQHpMsOHWzfvMRZnDheBb662zpxDZf
dQ4eaXEWuEqudk+3KLpq6oQxYf3mafZdF0Xr6fsYEZZwMmqEoAQNeDl1X1ilQfmo
XDJn6s0gJ7LhNduuUlnRhR1AxElFnGJQmL/joD7VOHA9WbTefVgXrx0gko3J1dVD
Aocnicrl7gyYWtSIPPgvYzmEkhM7NrmzRvdK5qK6swx6RX1d8Oq3HoX5Sq6GbNvl
ull6qKeK0vdzM66zKkrPMk+8nDe0NT6Jtw/sW+HMy3XKs5upL9hx5L/5OUgJkgdK
2eNrD2022v5aNbPJ8URu+FlRvsu6J0Oj+5qhwXBBUlyZWE9DxDonUJ7LnIeUqqmY
AtSXIywQfAEKnCtfNeJecHCEPokwEYmhTJWLYbM/VgdG3PiAvsjRwPjdFUc4Ek1x
20Du4jDYQPLDPVEapQ7/BnSwbmmnu2P3x4zEsbSQc/qjnoCAOzPk0QFAFDVHq3oI
B7aPdnq0I+ygc0pK6lIUGbqC1I4gQgzU+7CEzagph6X7tiVlBe0bgXUtEJo2qGzu
uAThLkxG/VUsRETF3oygSEdce+1RlxHX8hTFKyJYH9ltfLVtCzKBMiQfs8UwcGSk
LO445H6bXXG0Q9qoXF2PymO7EmPE5rFuuqlX2i+f59Oj/ricG048JhBvqOFGfc8q
tuRYlCiTDs4uoeMxUIxktut/T3UXw/7SNv2p3hWbghLF4SPjORVxduuzIQ3ehxvx
TYuklHgCvys+328Re8AKwc1kPAGxuzeb+ENfSM5y4qGrajwH0pQfB+rCa+jvJfJM
Crsiz4fNnIum9wRs6DI2eYM79ivV8yvRe96K9KGyYrbr8TPaOCwlUXQUw6JDfcbJ
JmJ7zd6LIlEn6g5bpCfUc4oH3wkKgO9V6r2pueytVsjwOL0RtN+uT9VTm2YJO1NA
iYrp5fFwX/GfamXaZ8nempWJcSU+nervrWtr6UPfznNIpB7rPr+dIl5rRmPd7Eiv
Qa3lgTkstANp2s28P5TyuUnldP4A8Ot8FMJCObeZpJpkwCSYJGzg9wgzMITA6khm
bhzxhTd6lgJFOgSWw20k80vuiRCdEYtTQuZKvtg25g4TrEVbGSx6k8BLl2JSDLok
Y22J7PEgh3Q9p9jBUpcPK36j4pZgZ/OXkNysizTEDVQI8Pf1vxKpR8ZSGIypDsUg
p6NhuXBReRMT+UZyz0y9rcoth59N2KTgagoAfQbuFUGUAkeDMabpVuymyOQBgdOa
XUnWlJEYG94jjiJYvQsWATs0iMWU4Cv+s2pnP/RgMucSqWFXbFKgnlHnBAWutCf8
6FZGPtguTR3O0BAt+CDvDtrYv5N7CyO/dYHMEfpQVqxQIX4a2rC8JcyiAVawfPsO
Di35wub3DJiQ0V46ytmCvfXxCUWZoxqypVbm5CI+D2TC8bDB73VdcxRv1yhyyxfk
WmrRuSwGXmy8TZBRfZx4YFdFCMFgaNfPfXmUYCQenQWXaNeCEImDtDh4rNUqV+dW
7y5BiDAv0H6Za48ya58nRtxP6XdfprJaKfkdEyipw85+zuPslV5bjHV0BicSfa6g
5ynwS+o5b5OUyeuVFlshA6aTFPKVt1Z6fyTzSmgmGCPxdEgePQfoORrCh+/3Gx8y
RT2/OXDZXSRSXipG8cp9uhdwATznemSSNpAvhGm8ROpaXmwdL8uCOqON8z9AlOjz
oBtw5CitF2eDIVOVJWOK4/Hkml7XBMDzO3LzRSzesevO1PfYSZVSJOf2A349ZF5k
wJjuIJoJHa5XkE97LC02pLKwwC2ntA623An1qd/mnUb/0TNn7dp9HYLU2YJY82ty
+roSW/zJvX4h6etnWDDrD0lxZ3MDRsJDkKogHxYwYK6MetSeeR3PLF+9Et3CiXzW
baDa27g8F8CYrhbYwI17rdNUFaPQAvfqX55ym7+SxPaKrfUhiIBmkpGlFcL/Yww1
pyErSU/OkSXRO8P9+JGhlwz6lm1yuXjE3gXNT6LuqfTCAb7R/kg1OmSeYO+cQMtc
UdGIDbTAuWOBAQdqqw8yLCWWe3v2eFryPiw1F+K2dKCrR0rmwr1UdVf2KuXokibw
D77zUnDIepvh0jTPWxmUns+YLJ4PVZosBk9BR57m0BwcdduGUiGqagLi+va5EGeO
o7S/wLJUGt0iMavY/A9aZIJt9imGI+9S6yJ56p9PzlRBDfe4KXg5vz+U0UJSNmdM
89uIMNiKc9m3Q5FXs38AVXnSQWxhUH2NyqRIbQyiqdevwcozKw0vWqkNwgf2N9oD
T1RPdUXEqmF3FJQorWGC/pd3jsEBUAIvtnTRMc9bNoX5+d7jD2sRTnrVn4QDfo1Z
zOjm+qDy4jDFSS/Z6X2N0cBL4UqzIX0zAFGe5QltURGA0Dg/lQ38hsucQmrgLELH
pc7QBzky9rcnXzJr81u8q6JF3fm9lJZAtplqXLNrFLwHOdHmuYc2UUb2rHqHy99w
wENQ0gsDOEOZzV9yimMfV712Z84wNfAatMusrselM9U9azak0vB2ntGs4YhInKvW
/QOPtUWOIfVqHJr9YPRBlhTzLii+OOI6SuVlzvDERLVxO+fpKCVkeLX8H/0UU+4V
tmFAQtlnH6CnvZ/z6xs5WMWMpE/9fbL7wDfO/lb7bphIw19+PS0v3DnRc6KIrDkv
NUtQsZRcJ0H1+F2C+QJzesreH0rLWbSn2YnmRSVxz/jkdyV9SM/CzyG5g4NTInyc
AHiyEv44iYQ18a6M3+vt5Y1hx8G5OXSbJl6T1wjL0R/+TliIZV7GXlxoWEX0jVXD
V/pDT/x8TFOeYd5pH7ke9/rhUzMcmVlwXo1SwI9EnKgMcwU9jJZWLDIPDo1Mev9K
05K3CbqGJ0GzVc6QsEiIyyOo+ugIjVisgEkLz9e0itb85ldmBmEm2mn7TuqvU203
EhuZbri+O2Hdhr4B9u2BucvkldZKY5kvjV37d2ejnMONYtssQSH8WF5LoD/X+Ys/
WktnW8zvnGDtPB4E0XhuSvMG/PwnoE3jwYfCDkuxqNYxtJ9oFkNoGg3i2yu7SJGp
cO/6k84bcprg1/4gZJ6ZDA/wn6hErR/Sr89GMKv81/Ackffl6ZfpJtx5ryqQOKDm
5hQMqySZriKyWnQqGqdrsBOJhYnJoFMYn/zZhUFxd4DJYEpdXsoqYYQ0csitMoC1
njLCc9BJdgRCZsLysU+dOVL9LtNRij0qQiLunNln50EV0B/b+gVRz+P4owEKrzgC
Hq+emH1zfeHVLcexY7310skDYZ3wlCpRp5Sl28i3eI/sb1D82gK1loCUPJeyYwWa
XGcrL1W+MVrbBHT6S3b2JAG+axq3ZvWMWE8/exggz4KjmR9nT56GgQ3rzOIQVceR
5phPc71/YqrfInR1lCLqLRMg1LFz3KjsCgv5BVKD/rnQLPKF87eZwmEjCChQ2CI4
di2inTacPQK5RDd5RxuIIZCuLpZ/05+P5AeTvLFk7MlDkjtArAvl9YcoMC+56J9D
doD8L30bNbhtvV8vt+8oUeceGcYdiVV6DJ2UePnajhID+P21mctudnhcB5J5Y37a
bRE8HQgo1gUfiOUHcWHd3u/DiGBLgc2ZF/EiscKQXIqwRWlTmxw26QIvP/bM/hse
Fp1AUMpuPx1FKJINH18tdIi4Ur1OOCIVQYpzJzdC03JspMwAOPWy/jvyvStpMTpj
eLst8pATxAZjGnGS5HxPdoS+8OJcMo62fU8+WYht/96NJpm6TdgBPeFkHaNQlboV
G2PAfECq43E8QwCO+RIiN65H70pqqNp8A3ea9zu9LhliNJCTEqbbH6k+VLpCEiyc
CHDZKK6GsXfBO2rQhGZq8kIEaVNs3+5ix0qCjbdW03xvywCMMfvYCRjvxcH5Ii+B
IHdGIbjdxEnw3Cl1wM1wSHGQ2DZr8u0OMU8P+u4sw/2dMfu++TnS9g/gIJoXFlVi
StqRBD8I4cQoDvNgHNwXDWMiFO4YwzgKm8riO8N/dm++VVRL/Ry54thnCKcvueCg
pYKKejLOXO7HY2losCcNRnZsjOp5sNvBuS5la2F107vg5BJz9lAXA84oyEIEh+Rx
12kLlDeE96kjipO7cS2audzHOA/v6q+hTFlqXuyrlxcNfhWN6ReDBTL8gYAuVDkf
FFchSh9Jye5CVCxhYvaiL+GF/Jl8UzD1719/r3BEoe4MWSpuAaeI/rpSGqP1dqJt
eMAG4dl6MyK3GpqolwyVJAoHnJ9u3f1FolseWf06wZBZIDfFPtcTNgX7FhpV3AkS
cGctJCSls8tsJr+7WOT7tkFrgOk/8OMSZ9k+Hw9DdbE1mlg9yTPxIiYY1sdwQOJg
lluiPRlR5nGFmfgiq/vAzuA3z/+Z3ggFvoQkQV0EO+MO2eUWQlzGoAu0SX3i/QYB
tdS6Q5h6YGvsWKefs6FbIFNhCPF5MTzgqhPuAgWxMMneSSJe8QBUqJRXgB95NPj/
1WCQJCDhtAMR6IVYGUBVZrNtEsdYKJtXPg7jKbvwHP4eGbAxRMm8BFkneoDLASC5
YNgCv2w4oJitzp3WbQHEvi8ykH5mhHE8gNFrbACWHgBa44GEm5MRydU6ONq84Faq
ugyuBTQHdC7hxs6neASPajnQCVErKvWRqTjbU4HRTy7OfEIu2RVJ+NdMJDBB2YKa
i5atpxeHj6ozrWWwihL7I9UNaSOLU5mBErnzv5WW2JO19+X0Y/vAFq00nwtCiDLc
TH14gC1YwmRqdVgDinegeFMCfsDc5JH8B9ZQ8ApFTzmuvVTJL7d1YSQmuOmFuAyR
rC7a7KijebHkN0u4cfs28jho2Q0TSQz4HxoAAiT/+sTNvTaRvc8UqRrIQiR/yMvD
/VY9YO0HrD/KvBS6sgG2BCuG6nQs7v2jcR/4msV8e/pAwZgy7mBudlhTGib5jTMw
V7BPUHqsNJKmumVNBbz9O8lJheeuWrc5Xo7uqwbx3NDdzzHOx5c/Lig6AkHPgZXH
diGxe6pXirt3GashqYHOWKSgAjS0C22+GROIwO8DeStUQZgOYcq5W1Iob6MBua6E
2nqf6TAxCNoRZVPbolw4rT9Q6P+GcKkKQs/By9izzWcVab14I8sKihLD7DbqvUt9
CsG6yy0b+Kxf+1+saeqJDvQQOIlcO1WStKqBzgRhDbj/ejezdToKowsDPyamErIP
XKkShRemlL9wbBfk3FVJc4gfsPVdGOcbxWruFRxXKanWz+GVU1WxD1ODk4b9yJQy
ViMmPS7bg1/Vo4PDcSQVt6DdmQbgN8XgfHjp966AQYINDZdLRI2jUTcNrJVYkv+H
phQ5R1VT6H73m0txhNkngAh19EeKa7Zx1M0TJmkQelLMiHzJtPBiqiYtH2tSwxy5
7gIJE9fXG6aJDkpVwcPOW70OPZsb0NU80kkljVoaEUYuUsA7mE7gls5pj1cXqe8v
Vmg8pPJC2ZJLLVKsubwOY1cVt0o6y8CvHuvPFLzjNeo8nlRrgOmiBC0Zhph7fuge
V7ozKqf80p6iaL9Gj7lOsZDD022I7HwwpNZEmstVX/OdhSpxYZA8lbzViQMU5ZjR
SGL6HG2Pp5WNN7Y+ZykVkAMODWxMozow0Lx388R5RnWlcEz5f0OtSuhwYvHCypya
v08MJNF2y6ltSF678PuGDbjdBCw0v2RzRgqPXGJk/ZMTCU0CIqTzS/xtm6koSdVO
wv/Dd1bQnAD7+ZAJ2HnaW7wQjGCBl4PBFmJ+h9NL6V2uljtqUx3t0yskPtKSSs1q
h0oWooE5VVdF0WLmPZmXFgZ81qnJGsel1wO3AcIfe0slZh/6gdRcnqVCDLpF532I
wHD3crtZIMup0C44LmYQhuRY4jxZvvN347aHpsTPgXExroJk+lv3B2/MEbVTeyin
O73PCRK8f9CRFSi3NFiJLAUDaP4Arn/pqyHHVZSCBPGdkeUOQyLUyLkXnI8k3xjO
a/Z3vHC6bd/9W2EsDg1XdAt5+0BsjxG0hBxtM5da6mHOxj+P8fnMOjFrHbUJSh5u
0Ss4RYYB6sUBu2nlOMHTbDkRZDCiatwcoi4StSeptCKkGiexBH9qLlkjSivZ6ZyY
CGkRlPNt7suDvS/pJECdMREA5yhj0C8CpnkUEREFQAUMrFPHWeWttwUuf85k9OWh
9XzD9cOiCK4teMGgugnqCXiJZ4kAKZ5qAyWjkha015xW5bgNNvLGcvUSxwtWoNuk
zagbIVPzmgXEtLA1ZDofBpTxIJ1OTtLKwK8G5u+oQDptRl8+YifdAeuMxZedkztx
4WwbkrZjyQqUSqEi80chU6u9GL9v9MO1ilDszB3Fgz8LE59i+68u53J/CEVZ+875
PpnDq1QIUF2VpS3UwkunfCUykdT1+Hekw68xVlMfHks9v418v+nxIwphJwURjDl8
kAnzwez1awrjF2gAx5ejXVfY6MyFlb4itwdd0y+sJu8l0WT0/dGL0e1zQL5Su0cQ
glC1O3GIK6j1fnFnkIOjGykM9ZqwKA5xP5ExlEbO6Z1eCZGhv/vbJziaDJjfgVLB
bx+FsOn1N1OpwPAhL5FKSFwK73tk3y7FQascr1Amrs7lgn24gtjt+OtOlwJUhqKr
BV2VBsltfBLXtSyIKGvQ/jBgeX4CEIGgYwQHxc9H3El1culM62l03Bww0GMzsG98
0RSxMdDenE5grQMA+tL+3u+g+LwAquEH78VuNJIW0xxdKicqbdUuMnMcL7NgyLo9
BOc245FdOP49tJMDtIX3gU13aopVVdDZhgcsH0Q0A60bmerBLezDHy7e5B+yyTKO
QxDqQMbVEvF3BDr8zufkRNognFJM14iyOA9yOe+uV4v2eKIGQL1E9TmJWxbzBoZF
Z6MEoNpFAt7wVzq+9op3ChVKGjpBNt/qs8kRhkuib7eBtNAvn5iNfCaD+fIUevgh
EIt1w8itnQpvqLhswNd6NcMHDCwiAh499+89kuFn26UGjtK8i2M5WA0QspsDddhm
fAfBg5+YjCCxeviIi64QA75MsVSV7AdNJohiChSnMWOQSNlK1AxAjTcTEdSpZ4j2
rM4XZylAf0bi7dLC93xAkccFt0XkIYiJALsRuCNqFn1D7stbzLk5FDw+Ui2lTO6M
glS6L99lsBTGGvEy+b6PtsZWSyJH5NU8A7Yhtk3pkmDHft02aXqx+DwvxaucDxtb
I6D2KGDTkBsFmhIShPUd+cq8xswsxxPxFko4mUo55jedTLWXmvKRKY9gDoW5vts1
I4eD8UmFnbdXJroNpYrAOlKPbbvgjmIW/XtDEZv91U71hocuD49RtAGZcWAfu1Ni
B8i5Wsr+VW04E31P/x0+zNuzJ0+JKcIrTGdGGDB+LKnL83+PZTuUzzdi/DyhldNa
hL6zS7euHwVTNEkBux0voaF68gruurRRRbDlLKMDxSJoyZ7NM/f0sQ8FGVC0vQDn
IJOFlS054p8yCd2vuFRyfRmfyWVzzgyyCxVa6cCf2TU7pKLqG62e0H2h3+H3odYW
kU4dK8c9AeNv4b70jBeM5dqK7uYl4dtEJU+um3sacdCc2I78M9ulVqoVG218bxxU
8d9XV8qu9MUY1aPLd5d08lVcd4Hg6o28dNw7Uf108dopbDAZGUpzS794avOfW1lq
AP7+Ij1ji9ON5f7ZdSC2t8zDlwC4DRkiiq7Q4DY8Y4A+nIvQc+6uxKw/8+LmogTL
cSHsSighYxi8Yt3rhILpCe7yO/n6UljZcrf+NONbMnBZxIWiasl3hsZREspkBg4H
8DRkIIiiCHGrafxbAXnLcxkzpcBTGkPzt5b4qOFGgi4pHWS+OwR4JhNl8x7sHhdn
+xMGlD9FebDQnvb/3IqJIWzBsmAYQgVu45eDhwpopk+1FjCxn9gafmFOcC151dl2
5Wz35PcNVmbjTX8E4exmDNe7dTrJfuQKeXTLOPWyyblcXk6qMIJ2912IEaQ5YnD3
PnjEQRE8CuPdPuvkyABYLU2vp3ZgzrupggmdzSYwaWQ1J4sf/8A8+XAVxSGonkqg
XMjucLwSW/SE42lrv+akqfap4DOrfKczIvS/iJLxDj380OBCLZod2A+Jx3B8uI9I
+8JlY5GqgdsoFdB3tv1TpAoiphScF1gWXmQ6znzTDT/bZkFSmx0JRJJ9xihSsWlW
gw8uLP5oHItA1u3/mbhWCatRFm7lh7RQwxrNJX54PpMKGMEWxRyFXmex+DReZN7m
LK0ef/ZkO7CZF6ffkg1aIb0SmP0xathVmXl7XtixWRGTh1SofB2kmMRqAHwhcJwE
vGa6xb11AsEDY16yQoZULGdXdGbqrdC8kY3LTa3/jB2Vj5xZ/YBp1UxZJv1T9M9a
b3qRM8n9aZTzBjE6XlAoOEyat7CH+QplGmOkjM/5PLlwZG/2HUlFz5JY2a2eTJ/0
FBUHjYHfSNiHtn2dMZ7q74XwmdWdCkELgsS6lyhZdGnpeLvJj5aK6XNQlIU8IqeD
WjDG9WrY/5dCP+4eZobbsY8NLUUkIMIqA7A5yjId9gaBSL+SRQ7zdrVwMziv0l8S
9ddjPWM+HWNTNXIxzeTqsvOHGVB3zMzocXl2QB079D4b5wbuBHsOcgGMJ4HO86G/
NEc8lFuFBNaz7HOPLdUdV5zuGexiOYW2bMnUjvpGVJzabTPyH8bHXKK1PwspCbFi
y3fKboHnX+4MhUcFpuSKpZ4XVMIm/vJQT13OnRDZmoRAkCgOBlDJ27ZbOac8EmyV
tWq5ENOAIgC178g/qR8NUhgkZ5e1fu8FWFApg8btGAPt0e4vbRri6aEDJuCJ2er/
exw4XOd0wAWoagoXciiJLKA3UgoH3cSYajGrZbC/r5jaSCK4hJ9ckbPqjSLf9l43
rRLFaemsMJd/goXIzfk7tro1VwqHENwL6RnKwiphpnAdtTS8nFLaSll2okb/FQJI
kYTNugE4sSGlY6m9SEcizrtmuUgJMNG4s/uKus5BdWSHneh2Vq2GY6zAexq38Ve4
uVgbn/jsfvL8OsiFOfOV28ec+EciFuihc1MLNuNpBdkiYS0naiilKGVOtuSg+fi2
eF6rHn4XtLvhD2R+jVlp64Sw/zLpgE3ySKFl+FhlQl99szTVOSNrbVR7pf2sBuul
3lbKRUk6vm8hL7Alp8ew5KX4RPR2z30AMYHDVG9BTNlFgEQjWSe60VeVNawn+1/9
4CzgbU53o2e/APH32zS8aiJ9IE+FwaesAdkDgc7+dB9S0kqCf3cmQAx4NLXSJY1r
gd8vPyd391JJQ8koJIxlTrvgO95eEX0jUk/EKCFggsVTQLFZpDtdEi9barrzA/LI
msPmI5MmNCyKFhbXCFc8H26Nzy72bXWraEr+TpInTSV2R5VHhPRJ3es5/p1BwGSi
SHsLiKfQexcDmjXNSmkjCWTdNeyf6r3VfGKqhcWj4GhEaRo13f5zco8K4Zy/Ucl7
mokqWjeBO5qczUU3NDxemi2ynRyf/apj7RiOZk5mSthorihnkiSx+nDhTnxJ3WhX
cadsi1deLlX/emQHb3tV0ESBaLgRb1aOKKvqGOAVD7eglByia/Y4LZxds3VJTzSo
I7mJtE6doGi9ZgH2ISbV3A4hp3ExBoAIMJwS6s0gv0wq+Jh4fdnSfdY839BAr0r6
fISQs2XPiqU3JaLjTzK+q6RxGH6emxO+Wb7IXn0SHvnuQW+DONEBS5GCCW4Huul7
hQxA/lEVBEjedEx4IX0Ga6FdINFG9HstmEPMuCN9HK+7QeWP8vNMkw3bY8tLUaek
TQmnTuUXtKc5GEGJpjSck32H2j7CB9SjmhKbhM/lt5PgEVQrSMldT9dkieFJMTc+
o3cUCQVA8Ii5PNREHIUmBC0wHIjkJGzVcTGVy9WqbalxEuq7A+inrKq0SsI/E1Cv
qyK07hMGwpkivzYdrSH54fs4SCS6QCMtjvTAixGGKlenlU3xLB+7ysZdVblOd7Bc
YY31g3BaUSm60HjSej97+ORkpOCw7Wt+0Q28MHV5GxbTgagThVSKiA04ahkUxRQM
xjhctnDo0LWsZc73bwWbd55Kil3vq3coUkLiBAMShFclEij2FJQk0MzYnMmGi3aC
eteW2DL2uCOArqfEMXffRRvPPNc51r0Jqy52Q7u33AE3xwItcfM7/dLTj7+JSAWG
f7u8qKkCrRdjHlnLheybi4auUCuq47ZH1lLLaQGGeDzU+uF5I8iS6444gk7+XDLH
Z9EeDuqz55rs99oiQqxZ6bMYGEJ/ZhwlkMbO0pKgHwKCraFWmkkoo1e/Lu5OhNEA
PMH5jPobE1kVArPBopNVtXMzyVAhsSZ2cluc0Vag0QxLZmE/VgboHO0tjVjVqDjY
6CFHdcw8a2TctuiqvzZ5g8CNCQAFZ4YJ1X1uODLnITsfrcz3NbTJEq0mYhQLCaoR
+FvtkmLYruSrDvaXQAR9XMVOZNocPWZN85J52vilGyaxBY2J1HD+9VVDCBv+zEU2
wShDnin1O78Bk5gL7kccCu3q37rOQFjyhjI3kIiWRhsYcKi8W+nh1ped6nU2lyNf
MFegQijBm2PMeZIvoN1BrRoSRPtaLFOj+lLiL2XtsQ4Kkc3Pr7Sgtg/2MfvzcDu9
vmQYuYUPwnSeJzKxJW31pl5trKGZhDHB8Z6aN1m1aw4hbgwFdiHfg7jJHPfrNCP1
LI9fXW17FreD6h7eOrY/zynallPCVyPm9c6c+VNnEraTfKPvuufmHT3tAmPd5TBh
HB1o0+V7XgxA4wa/X/vm+JbMFNDcZ43kiHzQiLKx1Z0ET1J7WhoubUtXW10tVSCS
KyGUvFDzzWGfhlG86MDz970DLST3+h0PgTM/nTUPQsOiTsX5n+25yDOjUfgKwy7X
PjHALXz09QRkT/1if+QtKpPy8Rm+M2jcZ2Ba+/OyWsIoYtM1tK0gYBhvCJ/gOVRr
hkAr0HEadey5LFaORLtYXWlXkkSKxJYxRWuOmtMHurzpGBaWGlaAodvmR0wUhiI2
oL5PHxdXw8ozduxDeQb1ZZKgkreradVu+snY44W10V92i53oFHZQM8OVLs/Pausf
EFtLGqKv2qSsCnUXLy68PkDi95mMsF6K0jWmDgcIMPFxOgoWO/+6bB1Bmribi5kc
ZzJmm0caPn8VfYcPS95DgWz65chbnleIdIzxT1Jr31ghXfno7DEjRrBZGtNIds13
uIEqVwgN5SZfyZVeimjp84sd7RwWfDqhtGV90PcoDsCIvkcKMOkHTgEq01mMAiiB
VTKgwd6noXiUFlfjGw5GDkqkpG4+hHhQGySUcf/Ujs1dAJhu5HePiNLWauwxHcYX
JcfuwDEOzNfr8xUolh6fJ1of6PDjfo4Ee6+KrRIQMAt/7rAJsg3lON6ixPsWpst8
biBvZPoy9gYf0aklxQ45IoQkTg5S8vtHAkpm2Ul82iGWnMtSO5GLylOWiGtRVeAK
S8/JAfuNPujgWzogRfYXQvlhORiLZEhnqCD158KqFZOXJZVyLN8m1mmH1lwxpaN8
D6gr6Hu/+4FtJdtMfqyxiqySsaWXZsus27hEib2BqQTHjtAlyBVVOlBEPnjoAKV5
bIk0kYpWnTr0ARbXV9POd+Wo8iw6X3e2oA2QM9Eg6Ih7q83yYZyVnaKKP9gpxjjJ
2St11g0+/neFu8zgvCR9k/NSbg3SRj12C1kTAIh3llTd6Y76N4rkQOkSp45fwBu8
A97KVzQjsrTeD8DvAel0B5RL4ChWunJsikckV9RcA9a+6w+vvWeDOqUtZcnmr8O7
1Ly106IRs2kcZw9Iii99UeqiY1rBpS5oZgH2HPiyi7LAa4DY+4ejL/f+Mqt4ysjm
DBPfm1ZVYXuO+e8z3RLGpsDcMiiOsvQJPU0KdIISu3ziZYJaxxb/5z+C29f0GQEY
6V8J68ndlvtz8E7QCO5Tvoff0Gi0WyfwDkoc5fQfA3ikOX4oCvWzC0ngfXm/YOSx
5xZCIASnwhL6x5CjxV2zo8OHlumeKJANosBRjXBEz4Rc9BctRCsmB0K29NswDONO
8DrEwTts8BCsQB3hFahq2EyULtIHZxSKjxUUjRC/Y18XGKFChVLKo/r1th0Su5+2
rOv1JHwWePvST0vWU9h78kAWE1CMCmB18F6dukzvAmAfrCxOfTdNiRBAJ9tgm4hm
QRLVrygXls5VLJ3Ig1XvjrxO6D6iZI5k7a2uwf6dxPpzyjsntH9wGn8AkakF0EdM
h9hSa0ZwxakVym0uxwkdWGzbcWFBZus2xQ1215S8UfezMGEDSXEezflPN/KvDRXy
C1qBRbtGjO2COJceDB81nCwelUhBS6CtUyaWHSXRg3ecVWGJY+t8qFdiYih4+epx
y1mI6ROmVwqFQeBg/Ml8vhltKddpqQzaObzRlv8RTwz+xWJWYrwymdQ5786uAOKN
3VRwnMCHkkrjte7YvQ72KqBgK8A1UbG2v0HG2t1wrMmI+XA/fj7vh1mA8BStOyGu
d+NiTdLa75h6KT26apvndB08m29OaoXEnQakZSwRpNrfsBXR77tMY9Kxaqg+Yx9Y
W5NBVpTF2ZRK44FSLtvwgMPGk2LZtYmspXf2h8sosjhJhzAGYnPSSHIPDdEbZ5du
OzOHF6AvRhoIPVynFBGzhWXd0THHPJFtWVlLj2P1aGpO9cHz3mv2ElcFObI582+4
OpZt9OYOPcPlFXT358JhwJ4RdVUb1zBgpA62eNzXGe88p+hkhrYo9YSy3d9L/84c
V4qzKCegcvWWI6h+t+hhmK1iTV1LDtu+zU4JjXTbNfp8nNAO0DZ2sf82YCzJ1n2i
bgBTI1kgYdGBv3vz9cM8DfS/AY975uSgcs5cCipI3PbqqZdaB4IhRgRYnIlp9kg6
suqJGWKWaKdy8cohVACK0qUsVuMBf34fHwGPFG1LQpGwQast3ZCqBwZ/RMnOjlSe
iOzWNmV+ZNXbYYSgVl1hatSCHi9g2QRFECt4jhs+wq7YH6RpbpPrkHHRilyfYqpD
WATWazGriB2Fj6b8q6tmDdHQF08cSEC4h70MkvpLigTnwqGdlHBfHalT1vAaCuQp
kqo/xtW+CratqZhO0xivS/2tZiAZtE8iciNWRCKCnrzzB4RSf5EMToBf9jXKdKu/
rspXLvm97GdD8sDH5POiyilwTMFqnWCmVEDxh7E+MEvarJWKRlfwkassxmYuCfeX
7jQ5naPwvPQkWmolZ5NyfdKu+qcZ/rX10OlvBrgtFY08HHg1tlwOpWalqcSFR2Cw
ZozIbqlrCaav9EeLL/u62RC3fX0Jw8UQHzXFIsg1byDxDyYaGGMrLHKHM9HSw0z9
M7YoZXXabo2KqSR20UpcRw2SRcLIrI19pwUxo2QWCIaIK1cnYFacfxVmgcJACJ35
LzSBFjNrqXYuTYRKkS7OUs5fm0We7ZxpyUulOseIbhZWxPpgdOxpbr5Awq7q2IXp
5tvRlyHgDbGy5pt60VJ1ipKdoYCPMQefY0cnrum08G+A2UTyhWsk7PFrpkd0FGlh
asjscDeKKv0OlmUxEwCWbj/8g6RBnz8teZ5KT+ct88aFlIGUDOqD5bleVAL4CmS+
A9O8bfx5rDKKHKj9oaHu0jp3iqdKlHZA6Q3BVBxndk5wedQBLeOWxu6tIH8ReVTe
C0zCx9qieJ7FdkVqyHEyyZQvPdQk8W0jWRhcktLo1Lb59PEhWvYkVhBzG5vxcA6n
jEyZqprauZ8svOPncay3bk5finp+m/HNajbKHNCYsx+FR8cNWWEFP7gvJhgK7Qs0
f4ITy1nBce6N/3svSly6nmVLkzQJnPL53HvTMO+PS8+2oVRkW4tu0+66z00eOd3c
+c4gxELEWuzW0XlStuUaJlMZK3Yzio5Q2wIJWL+PY6tKg/N27YJ2DD8G/+EPw4Hy
rD+KkAnV07S7YrTktv+zcrVCt82KHQgGFDPowx756pNHkl0xI5avKGb5sJzV4kTK
HbrECwHZkKrFmfxCVtxVYeMYbCpk6YU3c3n9xLsX6yZ6WbNuMftZFGpadHEOtT7+
jUCFzfW20kVEl7X68DpL3bAfa94/dGkBPBqn7rd5wh4gYvTvsCWQbp1Iwe/inPhM
FmE+NlHAy7xFx239pC3IoygoZCI7oN8io6t5MVA0dG6Rm3CDkS3rGBw7MLVBe1A9
FBQXctycHAjmtky+p3B5S4dqgBI4M2goWee90StfQ5fjhHrEZhxhddUyn8IO+Qzx
mpWNbTkUGaWuRMNLtfnGeIUvkrXnPrUC4Fa+yvjzMj4xfdspndhosFAtdkj1WWst
6RoRktMym6NV/xah89KPl1nGyaMu/tzBTjGpUtA0m/yQ8l8d0+xqgiGlWOvKIYPn
KLyjQmb/g9Vys+Uiz9Hqtr8zuUy6KQqbr5n2SuYWw2d1eqc6/IrvbDDu8obP+yTp
USOJXrHuFLPQZEMWbCar3w9jTo+CXe/HHndWXZBPLWpKThYdCheZufyWVOn5Yk6F
rhaUT7vjb51ZoAVUqnE6OSxXscJ10ie+sZeR65uibIMRdVpqJdKxobWtuZzvm9on
KtILtH8NHOn/akHnEULrwiQiDLaaDoanPUJyuRl0k8OJ4UW9lHQnUQ50A1Nb4F25
kXcb2tf/F7l3gi6n0kCrf5nADfLgNjK9M2SSJM0OF97JXASbnya9Z05dkEPY/zmX
aZDfYhN7AynbuqHTwH1NnkO0S/ZZjQ187gn6Yri8HJTml4AbWOTQ9JjJsM3hlfHp
ObEyplSYsvKnrd+1CunzEwTR4BN/8Jg7AKVjRgPSeGuVSloOuWrps4oc0aQ7cX0P
i+i36XxtuCyUgsYKYfTCmqf2uH9BA19VXGgHndMa1h8KNPsx0nwsSs8B6bNm5Rw3
amDHq8xGxM80wsTFPhl/sqk497kd505bln107e33DfLu8GnOa7nFl5/FHk2LXi6M
6uI7zjhAegLIx5eHbceSVN5IKKboW5LdX8xRixLsA+woS5pWrZLW2NkOtM6JqE77
ZKBxJhNKbHQyzPdOUbje+nRyGyrvny93bItnaYLTUFh7+dJUVs8LxbYOvkLOM/JS
NQ2D01B6qBo4oFxZ6fFd6+vMeUGE44CVgUFoD2nKH+aiW+eawVFJSzU90Xava4Pe
YuU9nREutrnAbGvftnt0+6vPtD5k0ub7UbfVN7TK+GAqrb9zYNJhw44hpmb6rn3R
vkvqVF5xOB02KHv5lDQDNzyBcakFiwICHS581L49cbaus34gaGQQqQE8gremdj64
bm7cI3lYoJkspvQXg6XPuKbdGsaYIYzJjq1wc5AuzPahgmLGPRO+j8nP7G79W7lU
Ts5AOMZSd+VEz7X9B1duB15M2cE9Dow2L6hxXG0633sTlVPPOSodv8CazPDFz94L
u/TrzSdUWg2d5jAiWDqeDocYbC/aaNwLzWP1m5nkKTogMy5s9JSGpYmRPdgKkSWi
x70bRJfhTuOxUTnnSlBNMe/vWBY41iaTsTmQ4lYKpmkoXc6J3ADqn73Uf08caL5G
E5ObPztShr+4IidgLidrPBX32zJLGdBfXftlNMZmZHyUJ9WySJJKYKm2gj4dyX99
34TTQWiQI46afFdUp9iTORjC4NBU1pXViLnjMJClBjbr+6WuF4aWRX7fgDIz5+TM
hxc041yO4rdvLdberONArqHLDKlrQf7yzRyvv1jNsM0fLQeVsx3J4s0DOVnFq2ZY
K86a2vVmcxoKsSWAn1F37mYbZeviM8wPgiCfPDq2B0xofLWEahfAJAhlcwuvp6A1
GtNopcvcbO4rMHJtPUOxBeER8CFYOecZI5Sn9TxpO1Mk50DwU1vhH/qzT74aQrWa
kTuXyY7dAk1K91SPJG2Hx6C/aRZHCX8eiYpW5B/iptztxozLS7gRFL4WHixDMzb+
H/xG/wPzAEcTFrJ2egRSA3zduJvi9xdQQOtfPL9FgzjHpkGIe08EM/GWICCx0Rrg
GjmDJYDCMsv4CVaRHretFmJK+Ly2MXaCsLZUcfrSkuW3zraTbLbLsWe/MhwBTyUZ
a2I+fNC4NMfSYp3+AfHN3qQ6/ZatFNtNpl89hWX0czbc3Z62WeGKVJSBtKKmFwMw
fcgXyO59GBag9MjZ8awV6TuxKRIJBD5+qaTCdS2TGD7spZ7JC3trNtNe86oMiSI+
PM0jSKjT7UgcZsV/JzHGySVYs1aPdlmx08Zml/967L+Y8vrViVL3sBUu3HfbPZsE
1Ti9S1pGTQnGEwt2gYyZs5sb2EK3jZyThY0Mwi3TJvQLtf1xGt/8k4e5LLlJYYUS
Qdaa0mevWqVFYtR3inOnlHotp/IfWYCKd/zADHl92vjF0MAf1uyBUa+6x9FPWTQ4
lymCiaeoHbgWQ46ORPqn+KzyCjvGyro9fyKfXCJUjd2EWPJ295d3Ixk7X8hhv4fm
mk5wQiig+ijSmeX4X3BQd5PcD/NSC6gXTiZFlrj5SYdbgoAuNkEEKnl0GqSeMlSA
5ny0qO03QLgv6wS8Ic0alZUvWKZQktAc0w4cfWRv0AqpNaAPl73yuQff58Dokpk6
v0zNHGVCrTrnzRXfJ5FKs/fTRg9Wtv+BLK6b4mP9wbeziCuF7Hh6JHQvEmVZU41Z
ZGilcWpimMa7doiJnb25MLcxiIocWCQREY2rL/iZbuyRs0gBOjiNy1u775v13C9S
O3knh9r/yIjb8PXK5v04M/uQieJCKTuQtjLNf0zvHAvqy5H91bES+8WOVD7GtS+8
9CVeb9dm4jDYn/JrVezZ1Z9hD72sLs7jBf2YWQDoWTEgF4agwDNOtOaldzGl5Fzz
E0rkgLOUJ9TQtDTjfKQEWi9LIGjvlfDmA7y5LyMLHRydCqDPp27ou99E8m5YAuCY
tHlxt6LkU1cM6u56qKoNjQJJa3+6b4LBjB+MuwqSb3DMSWyLZMyZst8ck+Fle8/Z
oO3zLo4v0m3sLCrCICROVinJ/HOI6shgz1O1/S/juAAvI8YTiUWlg1VA56DRxZE5
2i5y/fCZlZ/AZ8HkCIV33Qm0yCkbEqWYKxnjlSyP65f78UgaribteDUJl0iEHWc3
hS7L9dwJto167Z7zbmZZJToNxdTNS7fa3ngBJAegIE3mFJCBskOxZq2UUHsl2QKJ
8XwUIe7vpnagP4mT1ZxD0fgd4TaUMe/23O50j5omo3k/1aRuz3MOh7wOTiSDOlqO
Yz8Q7q5Dnb/MXlt/SkIloF46YWL/dqOlrrn/axM4J/04TnDDkxWaCoy1JnwCOsob
5XhnCnyeBmOCfMq7hgRMTQBJ9Y88UyAyq610G/nwOvDN72Xih+4HBHjDZcuIdgDB
rdthEzPe0+vYr881ry7Ann/PGZnrkIw6zAgQgtmq6fUJqKW7P4vKjI6Ue4KfrdS4
kw/N5xJER1DMv+Sgfar6yjBkzW6njIDDEHHJiqaC1xWtwKOl5tmC9Igk4yiiV4XB
MBHJI4DDq2iy1TPXErKDLhUbodyLjgx/MxRn4M9jJ55jNorczbC04ZmnVhbrm38q
oHggylb36sUC7NK305maUTbvojHBJZKvFtC67s6cqcagGcez4eA0b/ptm+HZwFZL
Zpb7MtwJPoXPgbXe/pun/MdlildQ0rG0tbLq08v+nFoJ3H2IFfNYYsFe+Xnu/pd+
Pv3x4LkIfnFiEs5hp4JNerjtY0CizMCWLm4MuCvjFyU16ebRN9JxFAylSVls9gsA
nVmosfbxK54vOylndW+WCSScAvTKxgL0n5vk//WlWLRWHEL0DEMj9AF2lSuHzNZJ
sYn22w+kb8rD3r1URsysOkBl6qiKdLIH8qfUrRDhoS9wzx8dRiaUPHSlbPwgJ5nB
MGS0vFDpJWN9slWRobs3RiVzFQ/ENl4RxzjQt0Kdlqzdv/+ALrz3Z+A3Iu0ZKzxw
W2r+TkWCbKMR//+1eBree4aHF8hzwTsS7D1u/vNuLqMUfsaUwJvsMMsm5sqeR4AT
ie3X0vpn3JVpJUos25XQUtF6lHeWj1sGg+6cRP5BanFvJYODHrBYhFKNLP1jTCyh
J7BtYF8dA1U3YErf3U5lat1j6rlRE6/LYBW87rt3dENNB0JJp3ecpoPHxzuMLLAO
FrE88kVffCg+kyFJXg6vmM4dUVSLhzmCxPIEBE+2iSToqfgkJTpMvzeIayI504Ms
04wzE7cbKVEpsfii+ihw3OmSO6f4ZwOZBWh47fvcK2qRhCJpxCGUwlnafQirl4Bf
9ZAAtwBjaBr90QiUspjPw7pxcVctBCiITjKgtpj8oAtuirfTxZb/zh8s72VwCHLo
0Drjo48FJ7oT1/LJr1eloIBlC4Rye8q/75Z8spB/RVVTM06vxHsVUZSjSWYvp4hW
R+gmVHlM1mzsYYVRZ+Zx7jreBEQ2DudxQkYvMDkrqU31Infu/5/JzL5z3kgvBvxy
lVfd6sdvZvTaRTZQepxvYAYWLHq6AVpCJZLqtl6uFAqHtabDhLUWqlYbD7rvsARF
3rTV8OQHUSxwyjeJzOtsK9L6h+SAB1odsj4+yMnzGBVz4jly263ZCagB3T+8puuQ
S9FC9YXob+uAUZptJrow7jMwR9DpT1t/2toQR33Yym6dDNdtFBEzoisCbyKNKidg
GLWeTL/al1D2IQu/WUaSExqOATQpTgWxO/qNJpgptslB7Tv5tYGBMhjZpqooWeKr
aHnm1sMATOk9qj7qGkPnuVhOknSVp4m4Xv7MjAlSbxgSxImemhmkqrbUtu0pvYs+
XpY/J6Rc4B7hOoACbGEjoqNGN6KBJbyd61fYZ26bRWBN6lo5RajQWv2rDNu1PTS3
YW4wQeosBtyU5lIcra22IqXBe4/NKNuXG2zxJEhsR9Q4r2bL6c+HCBqAAgn0Stht
6p2HpUoHX7FsqwPxyeQHDx4OVfo+N/LP+m15pmx5hFNl8Ad4pzF2PzPu8T8OR62+
evbFlQQF7shmTKeg/1CgswO4Z4/UkJIQQI48x5GNJCnwSaMDDK0V5g1q3vXvNt/c
DgLs46ZqljcMxKyMe75WE7gt2vYy1iErcc8wgK8qp3j2JVH28IJcZYI/ZoCKvlv/
73Y06Nz63m8OK6AxfRsffXC722uuYmxdH7Z6W4Wz8X8Q1zLwmC/CNluQGQWT+8Cz
DaMJpaVaE1wqNBLpwrXh4/LM5Rd/nJKcxhj5wGEWU5uh+JHhCtjBoBcAcpOUPhMf
cX1I60VczGXnKlRyA65HWgtrRJAFaLy20Pm6HKsTe8wTiKYh0lldVqpjkI9dL1H1
fPuuLZOjetIJ+LXk8LZPsnlrMM5tsIs5tynjVt8ZVIe+rQxsk8E5gJMOunCMb9Dq
S1dBykj7y9d0oPSV04J3HEy37UCdoNAMhvS/49gQWFX/Gzo1tTTkQsmFykjB+gE6
GMwfAHMacxhJ0T1CCAY+b9HefxDHdo0LoZDcXH+KfzN5zEwjZiiHDF5w7m7V0Laq
StkII8CG2DxgNh5PUKSYlUs+QWoPo1vUhon8gRGeMOrlideKSIc9J9EZ/ZDVRwUT
XDKAQpqkF0uNQa9zhIb8JXnW9FzPes/7kYdUBYOvaY0IEJM9/i6vqs+MN7vhCnjJ
2cJ+WInthzA8VtJc3PscaC9TWfMiCW2+zJPgxzLWeTSSswzezjCcgYKCjvf1Owdl
SiGExrDn0fymrr+RKIzONen+I4BkzcOK+Edi6tI5LMBnL842453a8LaV0nGRjMHk
SAHW6NC573Wjv+pM7yDg3vJ+0Ivy4fl3T9Y9IpffeIwWdMD1KT5xdmDsLQj15BbD
4K+JT5MAP9q4jB5+NbLm0h+BFG6nRFo+mj98FR3/G1MUz8Jpm/8FaZ+lHPQx24PA
S+urRkaxRWbBHpCq3UmhtGM/aVvb0GFq9n0OMySKbWRzjE/0UbEfnhjYfkuteSrI
c306JE78s5kbEC+wTi5kdtR2rVeCqKc8N37wArcyEcyfshjbu0wk/5U+FzPD6XrC
KMCtxXTtqsY7e0wTi0xHdoNd7xXmfzfZ0wdKUGdBXQFi4++h0NBzr4HmtY/85Cqs
7TmAIZwmejkUkmGbPRYCmnKBJheSVGX5RipleIeNX2/XwysvX12GCNdAFcimptMI
2neO4JtthBWtLNUzWIApY1V0NGd4MK+zx7sM0DBpJV3YlJ++mF/dm2elZj5dh2+h
MWRo92LJguoSG6qDljP/ODU1xxtMRDWt95PjrjMDahkv1DEYduGgkeowrCVE3GJW
VV34VMO4/iKPsrVyoDJj+G9ufeTWL6anqPDi1K+/mFub38lW+OQobfcyRq0TFrFf
aFN60zs0hh0EM47sAlk7j390/0R4z8QU4jHIyYmvtwD2609EpXmUfKfRScBrR83P
EMIezh9VgAgBXbRorxQoHv7yuDvUCvi+E51qboH5qWtazuybQyaU/uYWVMpsG/jn
BPjZm85OZ3jIHB5kA4jm48Th+/UBpqqkK72oOpnyHGkt2UKJkM4/sjkrZ+namacH
jVO4vorpLL8TbrJUVif7qPiEARF+mj4rxadJegjKXNvNdCgSANNi9xSz/D5cjJ0B
+R62935FPXHY2AzUFDq61RJ0N9M+/rwyA8vympTbTtGD/qdH7OnU/zqKVT0Cz9KE
MatIyYKej6iEMNmVRYxrl+TyJVYFgqziioSx5O9QiMuwBsBFP1qVDYwaXHhgpfUg
K/GmGhcpRQyTzQHpg5plEJ1B+TGHTk1HakTmxVSgyry4+k0G1aRSSUBgHbfEA4uY
UogcnHKGd1j/zLGoeTxHXHvD5CV9mJdV+tGCzPtHwLrZ+jOCiU97dQmYTJrymwbD
60rS+1//v401XDyFcw7iP187nZ/JSWkV91T4ZHFRv2MUsP8umRvn33FFT/4zIqEe
HCxPbqUWAg5EU796JI1F6CMKcf/jOmyr/d8RBh46B6XcVwExJ1zog/CW+zeOvh7c
nYnqoAQD7EZqhoAcSpj35zvuowvAU8ZYmgUzlmxvFzE56YM2IWS3qeZAqfQNbtP5
HyUkeSY9Xae/3R5XcrW11X4sZv6EkR51DgDBO9hfLPTyA6GvbqjgBUk9ZI/KIMzO
AW4fzmabuPT9JXf8ygDaqrwHGrOOxZd6rN16XvJDRzRu3XnJAa3JXLW7389t2iCx
Ro99XPGM33bMFigU/lcm69NwgyLWT2Ak3XVrJtMI/hXKYHAYXpAj8oszZt78gTd3
xMwAMrcP1OnZLCiXciHyKG3X4FwjdCxlzEttPURgzTA/jyU4MBsMzIRc8wdh1nFM
GFKu71OC772cBgR2LbL9F8gyzvps7Dzn2y7TqjMHYHjQWSwrjVsMK3Vz8pExTM3L
If70bEiuEJ5yvg/1FlopsWqr0YbF6C64SS7P8b8c6nuBbDW5RSp2l9vFxLt7kC86
gyok23PQnLo5nFk9iG81dAt9wn7DnDfnd+9MhENjxEy3bNEop5TdAb6TtazGZcXG
X7ekak/ZzTctQVAAhnRwBjNbr9TCVjvrlTcxQaA85s7+oj1v7ALMZHdrdPdm2JZi
OeTV6508QIN8Jspk4c28dDgvhsbQKVZevThLsgZq5V7jiLsERUgvxXgoka3eDEo3
vGSrm5PYXSJuW0W4Uawat2ZdQq9pfAG+9a+KJdrGltr6PWoQJYKqsGxBgorEzt7+
tS5nTAHjfdn8xkS+UpJXEBDjdUKwHXg2kj9zHZKN1jaKsqmT64PbDEvuY1iIfz7z
YiuaWUfM3sW8AQIBR/9qpSxbJ9UpuzZTERbwkY/jhi3wYvQ5xQQ/VeJKc14mndRO
PLZYI3pdwSlytFAnFQsYm29k51ZzEo5z0Ua7AE1GexrSv1nTqB0ETS4cE/KSgP05
qar2geR6v4GZFiTIUMJRN4m8M0xNV3PlukUcOW/v+uupMeL6iEnNN7IipHPxzCw/
JrxweoVAQPRj1a31YKrsZ3AA1rr+jLRqwbC2fdOIWTsYcAWgP2tO+WzJVWyJoo1h
68yuYNilz2+ssBTdb/gMhG99Iy49o3PZML0t+Uq/YFrmgRcqicCw8ptjnmVL0Y/A
+AXMbUW5F9DySNnmSseJSzt3xLNxi23xGYuUCoaoNXTu3CIuod47NFnBeHltv87w
0wMFZLPGa6v6Y8GB0iiYhK9VY4EjfYbO/cnhjnN7vBDj6cqZYLDkr4XZrpa+0VZC
/OZOsrSJ5u1br6JdL5Ctmw+YOWHjLs0Bx+XIAVZRY1xnEtWadpdGtOFP+M0bFe6p
7UFeAriTqL6xp3DEe034Pb7nqAtZIwsHSsh+pX3sKYhoM/FHE42w+v40fPWqW+20
ko17ASQFC5clyTX7ucLhvewDFaRoCLP6f8zOfwgBs86HK3gTNc7BEldQ5C0g4fB/
JSzjRFDGi9V5H7GzwstWIpHeg7gNq7viJ++nstsNSGyGcwxxTKH8g0yyYxOssBJn
k3qHfh+yauqQk0kpwlgXSPXkJYvodyENR9z9jazrpE26CcD3LVIsogKgP5oeBxJ6
9+A5tI9gDvWhNdUQRC9S6Tr+brXtNzXD/yBKj7sRvvA236XoOwAt2XE0WlWudiUO
5rZZzzc8xQ2YlkDbT5/hdxcprSyX/067lGbs8IDMrYQpVXZFRIXy6rYWawV6qSIf
EmbSGjE3Ji+ZmORX3m9flnRzUEqfUNBzVW9Nu86Hucs83CgxOsdr5YH0TydV68NE
1j8GWGpV8pBVzunQOX+M9q6EcKc38KFEmvNrPyrUhNKZ6WL1VccO2syDzDBBKTZE
Ro4UULsn+hEIEAsaTo3o9JaZbNDJtI/x+kDLiFxGIHoMTNPGJx9PN3+XXLipw34Y
iuyge4UjOR50oduCpkXjLdYUo3HD6eviRMrfQD/5vaZESRWIrE79LxDC5c6Lx1pO
LMfLOxUz1prPIpDcxw8cxkQrvokyYJcIL407lAW/U5v5m52CWXzDunkwnUZhDhGr
My93bt6haTUJWpyk/a1rhr03glQ8wdBfgoSwsbILsj4yShMgSDf2itfsjNlFMLbB
iVVpt9koAAodk86OEPjuOSWfddrrfzWJHT+q8qf8yOuwrUQBQGWoln93GP7Df6Q1
ZMhdZU5GeaMp950x7/DmovEpEoXnZpXV9LUK4fltAzivlj3peBz7rhhQcZt2i3rW
AqnrXBY8wdCHrXMZ/zkRpVTDAtNkx3EqLIpbh2LZn+IidvjDmh+Y+adHSB8USGDz
VXCUJ5rsq+x3nOQlx9QgUrCI253CVGWpR38We/ZWz7mhuMeEsyX/Fw1c+wv/MF4n
5unyXwcfIzu1Q2g7pq4FbZZnrBR0/BE+a2ogj/RYUvFT9uy40uAYVFjILQQDkUhx
Si/XXJOoAm7fLGuLR85hF1w/Csev+HFegmn2Xf4MPygH0NsZVaB88iQdzNbqrs+X
MeuhHIKE1DQGKsN8rI/ZycCGvW5BLDAheyCdie/TTscAh0kAvNU7P0aX0itX0BI8
HYbEjdu1xcKyuv/sc4xHvpp4tw1DToSE5sXma1USdfzkWENE+AidYR1Z7OAoFtG6
7jENO4fSlMnWIxAKw+ShWaIznO81YGy45sir7o1Mu01APLMm81fippizMBCkrjT1
usiJuwqfPqW3m6kMZMH3PXa5TTH8O2YIp0do2oExo4EFvDlpWPXfyK4s7YG44zCG
uB/bVPKy9BtKme0zPobPrTwwTgHnMbecD6aMfZ8O8KRzpiI0jMm8Xcih1/YKBqX6
HDlMaF9jV1KGXpi2dXcThXzNGOhJFyF4CqQ3BgUorc6Yolh1hNjg2RnKigoaydth
8/vHXmyf7HnIa6fZmraMTGp5LwH5TUuFFiM4YQNQBbRBwH8l+OJlbMA975CR2vyb
6xENUTa9nxY2JCHxWfG+ThvgJbYEtWAvQfBzzSdbnLtD5q0c/NJ0T7wD5r814vx7
v5syqFfg4s/Aer6Tx2irg1rmVBgwXPlm5jS5dbMgHKCySm4EAT8DLRmxVtXbcAAn
Qh0FDGZMqNptAFWVbTv3xYgLa3IQa2KzgATMW7LEu8688kVW4pVM4oZI0prighCL
mqYwWHy1yqhKrTAgaK7KhtUTknNS0QX+JuWAloVgNSSC+ghWLP4rlElFVlRLqrpn
aTW3WZ64Atk+DCY7cE5w5YgMrp/6MRUL94g123AcQ3EY02XAxT9wT6G3k5LT7DCm
WnoBWrnGZkU+GXk+vdjwXTA72nT/GAj+WaNyb5T88fAC4LY3wf+DMTDXspx/Jd6C
Y1QLB0AE8+5v6IRaxVtG+S8cdxPt5EyRHEKM4Nhu1a22SHwU2zcU1QGl5sP76f65
MoLAWbqMvXr4CjguXuGix+yPCsqHKuhUvzQB9mTzM/xxzJUsAviQKrdQgxZWELe8
GYBAWzrGO0AGOiiTHJ+1YFgBYj8Sbm3zjn+KO9F51dRV7BHzcNbsC20ENsm5FJjn
kXsnthtLRWhnR4tMyfHcpI9zvTQQbkEuTvybre4bABhMR7wwafo+CbDJf2lCQeX3
ziF0JIWt5AC14/fRcPyB8WQFt2qlM4KM+Fjd+/on9oKeLtdaoPN4VEw5/uMO4yy9
qbe1oePLyI/0iH09rM+23CgyE3QiH6Wq3bykGcyhXOxFUtV24e6lUtJhvj3yP6g5
IN1RB7aN1s3YI1RQwewNxwfv4DSoLemXa8TmZet2YRnRJ06Ym4aaARwFHxSYNxd+
dk4IXI2/N/f1+JAG8+/k5upkvQoyXF7wM3I91bae0tkOwSSW2iANi0yNHUU1VsEt
tEd4kDlE/K59WUpzYYuOTkRoiEn2VbRW7qJ90AYsEAA8MSeGgR28cKIhGdzA/pZ3
OwxTyGyusQfwCx8oWqlvyjlfejicvK0EquuJodEq4AVxS0cAZCemxljRIgui+h0R
F1ijvCqw1EDU1hq86yYFXoQ8J7wTbof5GSW8Kmw4mLVg6cKXmmlNDX89HSNNpxaT
zz7HURkgTEcj5xRkFH4d4yWPfe83OKc3vK1qp8DztFML9OxuqRF6hJCTTjRQzuJT
igbPGcbngzfWtr22nVkVyjGo46jM3Q60wdEUz15ycqxlDZEcmCmlJmGoYNKGZmK4
F4BYMCoL0UCZN+JQB4+xjuvDXhG7lUsI74qKWhGGgOYv2ZRfgdkOynZygX5QrHZ3
AXwVT/z3u++GottNvA8CoxBY5JXT112129Y+nu4YYUmEr0unbye+lBi8ctNbq9Qa
DviqIOmpZiTvMZCjuNejsXpuTC9432AXpBvlYCuFAfQSvkZvMTdSjnNoH7CW8fUU
yK3jsq2nVgqQ82hWfoZ4NdDGIwLqURFvkdDHUKC8M6BZ+UguQlxQd4VfSRaIgVYQ
rvfIAaHJCvxlamuUYTs7SO5HNd1/2c6fa1Yyb9oCk78vtV8IBgfrMHaq2ZdgCkL5
JyMZwDNW74U3c8dQDl1ULuE9NAyM9Eh/V2lEdmg7xyFc6fXncWKWFvxm/K82sO+a
YGN9U6m82ScBYvy1E5KDopt7AzR/Y9VVuGazsJZSpSpT+Kf+HiWvrRsFzqPTJuDM
pBOCdI6earaw2fyvlpkisrDoqe6JtIvEIiKw9Rc1fns/LVDXBEEBHeUxjmJg2xN/
nCJpH3NdLS50OaYW3k2A9xxGzfYpL8/ETMQgU1/5iPyMGSuDx6y3G+BQGbSWkZ2o
yfLnOc8f10BRW8aEZQBOH5L6oi9t9HjlcK6dTxV/tVwe8tOdZoFbJ/aJV+E4TWxa
YCS2iGm230i0S/3zw8kpd64XNqSrieOx4r83DzHY/Se+Jq+QDd5Ihl2st04HcLev
mzFHkp/yPKuR2d5Ak60ZMdNnKUefVlf1xQbudmvqTMeDxNS+j/Svv0EbAATq9Z1S
Rk9J4W1OKfgNZbDZK1lLo54hpFVTz4X0Vp0EhG830kbG/ATBr5I0+3141vjl+XZj
Y+x8scPndwM6e6aSIeXCwjANbvS8vUNkDjP8b6Fk+w2uPvnqQnF/Rvoo4o52aR74
s/hjqKTugAjV1YXIAsCGtR9OgS3BWbCwxWW1nnp1lvsyua1DaLWvIaUwT9UrT4P7
eytqsIEtsxV+86GpDj+2rBmwrJ1Zen8PYqcFKexjExXzS5l98nAJcZwt0A9Lbs/V
6WkBxWWiZQihPR1MYql3l5ShTgtL6+a6bpmpCqpEsS+xmhzVe2O74060aVxGs7M/
7SQFnooA54AgU/5u2QB2qyFnGF8t3phXYhxmGp0qRTWz07Ymhsaj993zMAD9lahL
In5RWI3RqwqvdxBp8PewqkwCXlqqMavogxtGpeyXafadoWnhY8+Rhg4HHKRwmj9h
z0J7bMJkD86kVgfTIPRfAhljczSdz8qgQmkcp/szkd3KN12I+W9PpKtgzQ+qaFAf
dsfj1bC3jGvOdnMjqC7hmV0DKNAoAH0P0LzxT5lsnjk4ol+hkHir35DgdqWsRqEZ
IT0YJYM8CSaZS8m/+dube41lLqiLs+vNUNItxrRoVAf+SIJd5wksZE0eXz1pfHfA
OLEdePA/ZvGxWg7mFAE3lw0wktDRjWVnAzZ4D4W0JWeM/iw/O4gyLg3ZYhkWuvhI
9reo+F8qp5vxftLoO2il9R5soQuYa9dDkWPXxYvPRSJ/my1w42a3rlZE1NoV2+Ae
C9HO6KDm9dl8fWPKTOhbRUwjRvjYDIsRHS/veTRrY81BXX1PVekptCZjTOohvzJt
cRshGTVK638G4jtfw9uJ9kYnShacgmwYT5+s/hhcLiH5o5AyT8b1eITReLWMv4KH
lOZhdyeVuxiCcqxLD2CXW60tWbGVbKlGxpzsKBeDzXyFm7ovDsVi+ZQWyF8muNgk
kTZ6rMYDG1YwHZiUqjQVArpwsYa6O9Pq0w1JT/T8dafNhSOn5uv+PtlrCrt44BPl
b0aM2Nrynp1y1FAcKtBL3WsTlbKm5ydVyOM2/Sakq1ZfI3DfbBBBnhCNpQPBRrVR
c1IFzk5N00M9AYll8kxVGnHe6Sa+Ki26vnaOkbpOmlMnczZw8dwODDOSA5a/axB/
6FCCuFDp0AgrOXJ4WzcSK3w9AV1HmSGHvJ+bR9l7IDawEofDTmr9x2FJS3CHr6Yy
hlsMNPxdhjgm27ebWnJ8UzafNBJo0gMApFNGSjnMENL9IBdALWVRLVDU4kKqBEm9
C2BU/9SzEtIOo0fdRDEJmQgj6z1FtzbUviKIBqRK91HjC3NZ6v3JYA0LlKN71tp1
12vFqLxtOmg1tIrRGUOacSTCqHtaUlfIJJjm9JYB9HBAUqUySVEOTZfGMLqqAQuQ
/9C8D4kiQqa2OZP0OSsuO4vqL29tCcT6wCr3EXi1KbRmSYzXOf8sytB1dhA6cWpd
9+BzI0vVdEmmJ1pJ3UK+IGTLQd7CSyI1wABnCLqE1ekt8LpFK9MhkyAHksw5nPC1
ikxSfqWckYp4/PYvJtchOGV/hRnXAXRFjK9hzf4L2IIaZkEvJAhbh+/dmLzL388l
qmyLJc8PXKK8gOC5J2HPNiBimfW/zA6+/+B8wghv5/x+Y382HPcYoQGmnI08+f6f
Legaa6uOHToEasXSbyG9fJ/kL6CaOIvVkyLu3xWY9RAlTK/PHeXeLZo5sbjqOtyY
PAIvtIShz7LX7qBmW/Anf5AQ+/eSqTK1r1mLwN2Q1sVnPhYpKWxTW9JAy610/f8s
9TI2cx7jkz011UowV6hspkzAZKXicuMpHM/wS7AILBVd8ry6qrpTXSKAaWPDVo1J
YcYX5QmVBXN4O9Lcj9HRNU3w8G/zfAHghgny12staZ1ESA5OhIpUxo3MyFluNB+w
UV6y3H6hz6DPFY8RUdI1PzM7uV50+qlohEtcnU82jrrZXpTUOQEou9NyiWKFJvzj
bFIOF9QR1DulVfpn2JML5nERfP4GK/keIejR6V42bmqM9vRaxzTbvZRroke7EmX8
0MkUNazgFzxaxAWZZFeo07Iic8dxHRbJXusLATx9L+y9ZMky8t1dZG3cFWn/r+61
E/a6kLULi9cJYBDT1cuEOO+jS3/vltnSipf+34tt9lO8UpsrLuXRVCJZp3/smlgW
fbgVbsIjW+BwmAJUKslPuVD1QTKXVUHy4OI1mTuJDAJWCk+bCrgZvWYRWe++gcsV
ePuJNFI+5rONYzcPWfW5+H3ozxehyE8D+nz2XiK4bd36d/48jsf06eQi6pmP3HYH
nrlta6i0lFmnHqx/A9CzVOa9zHzlRKKPjKVM/DCzoqQnCuEcCAoLT8GvmlVDm/+4
nCYtokGFDLYp17clfcdSJ6Sy25IiwxaYvCjcluL0gFuuBYXW3ALEue6BHspdGH13
wEkfzQEyNL72loxW2nBBB8OMmnMcEAcx1wP6H6Zu5tN60TN3pmP8lSYpNRvb3SNL
KCw3jmNa2DdosZKUxsze3AdeDXii+Y9UftK8Bv+SrsJ4IbPK402XdA6kpuSMWbQn
G8oNUUfAW43ng2jBp/z3yyTBTp0rG3seL4JaZis2EbvoFxERQ7+HXAyBwAcLJHtY
RXXBSoRCZvxZMdKIOI6kxsepUB78uJHr8nhYDWsZsunb9rr/kj1l/5Bzv1qmZ2ub
3D5LUaHo7oWbYQj1bzxU8MUtzeALmkbAGrPY3NWqc3aGEP7XpygXj2cSiLLvuLFn
/O/th3IYCYBqkLKT9Og7p++K3kZ5HHOEhHrY+zzoNfaorpY223k0tLfL0hRldbLt
uZblWaXSedEbf/Dy6+UoelK/sMgGMh+wkqBMe9QuBx+nFO2ZrkNHIqj2rWvWcvDT
VUPY5rZUqGMA9QtCdhWDfGvwI7skW6FqckZl3tu1UJ+2TzZ0syoQ3QPW0gzdzbSm
GbnwS4KPMd4Iv/yULNvFNG9OPjM8YZW2hzFmGHGfhsGw8D/gHvhGkR9ITb4bUyDn
/5zIgvxk9fUdzWv5SRG4CVKDGsj1rm0hmej6ER8fMMrOileEVpDkUL88pdmlBLwa
EoTlWyLMat8WY+bzSnu2kTXgR7wuwOfADuE2JWBEN+z4flbfeY0hq8iYPfQs1r9S
8mXU7Pg6+wK0VwHM/XR+CPp8kFA7OWkkfPeS8nTeK4bRB91zpitFxa/0Tir83ysJ
R+2PeB9I1gu6v3Z90DIMcSMrZ0NNNHmP5UfWr+C2i/AiPJC7nzjHcvpLGHnUiZ83
0iGrOXe2WSyLfiLaNLvt9ckZbWcVOWA6n7SZ2CdVp3tlwXU1OItDND4g7YjRBGVn
GQ0cqXW0bEfrQHwGNWQqtkCgAuusjI4GKSTJWdHiY6I6Hnf5OowxRsqw3Rr7h0x6
zsrQwG+qUTmnh4vfe1/y13i0blwnRy4e0rmyS8qXuDrkJekEPzrHcs8d9Z5XDZxg
WHn8UJDE3+95JLiD8IfbchCxlXxFewalanXSdC4KlzSoWPSk6U+JEmj0jabEDPbR
tjHhiIwWMq1q97PV5Gkdw+WAiTevkQEOIdw6DToXyyy43YN0l7SoeHKBgxGgJK7/
whKUCqAnbZKz5NkJ69C8zINMSYwaAqnc4pDZ+jvV/ejJcgVdiAUJ6VKYTj7QMvhz
YIw5DG+yqKReJXU17QFYnBnkLd7c2SxvggWxQ4qe209RelDPYSnOvA+hZKtEREix
Xhvk417P/zOXkXTXCSrRzCmuR0KYKhxJcaSA+13Gpd61efQwL5px+QpF2o2pjXMQ
+Oauxglqv6M/zrzVBAdGalGD6Nm3BIzstoI6rouL5fz7TaqVB0EqEBvUmGTLYEq9
MY0klMLAJ0DLcyzeWdN/8xErcMVdnyGSlnvK7MpEuAXcu4Ql/oxprWQGwkI+8VEf
pVB3NZqpBTJqxly6X4pB9YN/IRNE+ojwqfVjLyJGi3RYiI1T//drigqt8cRtzazW
HQwwWionW5SnTTYYUkR99i6SUmntX2e8xMrRaSkoGVwLrsBKchydMlyw94weV0WV
+dKi8WtUA1Ha6i6qiAJMK29FPrENuSfO9DhJnoLvn/RyfV41JaSQUgdexbDdaaZF
9RXyyfOGWcxjxtj/MMaoVyxVx7mmEYDev1T0erqw0QBrhSdRe6Ka6YmfT0a3HF0y
6cE4DeXPqtdLr0uwxd45BfBAeWe3eem2iwwEkOB0Y2Z2HVkNKTHBn65E3H+BPR9K
lDQd47wW7yjCTgvfnIUtfjscShCmTsltouHPR40QC5Ln6jk1DxcsLQjVKK708mYg
zf7WyhpzeVwC8kR4jMbuIfIjuVeiVaUz37kIPONWY3ncDXmL1fN40LFM0zvmSNz+
PF2L98On5CajvJue8KPBck3LDr9e6Np4iA0rcMUs8tr2uiNbev54RWpET7LeutIu
jZgdXDvxY5Jmwc54nZ+WNZx4ELL1xGs86znh37J9+YAnxKYpNK3+wtzfoJ79riAP
GVacq2j2XLKWJkr7KUYAeoKDSj9G7QRjI75dOWvROft4MLCwvXkzluPg7KZv4VXU
i47F6zWut5REPVL1a8oWh6V5YOFgJUyKc7h8xH5BINKc9vYq9Ryj78OWAK8S0ho5
jncD22r9vFA4nBcgUOWguhI2O8nIvA9N1PCMHDBZhMe7Fnqu2fvlYpht9XQvne6s
JvgNIWZBM+oYjfJtDeBakjSSNbe10lqc3q6tAv0oCaZvc5yFo85dhblYAXXp3PYS
XGBFMz4IWDO3GZ8wSJGxb4FyvRu8qtc4591xOrl/G6crbywiLU8qqg9vm6pF2tQ0
2b3yrYeZ/6wqZgs1ErS3TUVfESpfSREiMH748wkmBt+6SjKXWolf/hIORvIdkAS0
uFVUUtDiWL+kIMELhEZAnKoRBRP//mM0SlKoiTZqXhhyKzod5PXYFtUzjiIHNI2u
U175F7rCfMQGov995d+hbM1OlVH2stzSB2ArHV5XmBZUBDJNFVxA/aLvNK4aBvHY
R5GkfhR3PDnD2mbaVWdR/C4zVPoUThxE3zZe/5WobJNmzerUSP0OxZ8ItPd+RnhU
joXOJkfuPXZmvhfeY2pFlel2bapVN073/N5l6tTiZynsRgGfpivZkF2tUfkdJT9m
gZNtwfuT37htnoD31pLDAHYD0OL7/3gDx4g1bjNlA+ot5suu4QMUcDP8CsNS7eZY
LG/WbjuxPLaFEQf6Iqbm60PZITZO3jrlWkXD/ul+QYj91EmE+u+bp9ACwjePjU+3
VQ01Ggez9CcVnTo5fQXOB+KAyPd67pAevwd2tiog9/sfEpjZgwNqLX3q+3X32X52
76ujjsBDan3XEgNNQO5Rt4cWq2uU2fGSJEwEYB6jcqpusMWidip1dt+hB1V922NL
T7eih/rYg8lLpfKCuMNHTAtdh0MMq8/D6UEIz6SVKXOL+asn+EAD9a3KUuLNSA+x
Lek+olk4/4MnOd/i8r9ccMknH2P8nTkdz2XMudcAWYib13XVTqbomqXKuUSfP3A9
yeLtc6cytMYud0aVWzlbPOyFkdnYhJHhW5tVHdjArYjentgQFLwG6sQFOJS+cFQO
mGTPsECGpU767lWK+CnW9X+2pY0fL9N+0IFUHATiSv6/GOD2yfk8ZXokKv9ZAgai
4TBDMKGiZPA4W/pQVBgvJpO2mlHGan30a1gTv7YNsPCPCfFesvaVuPSVpOu3UvEg
RfhvfwuNp1v8xLG1uiCrDfH7KzuIC02W3ne2ZqgCpuw/gbucvKn5uI3OSFZuB4Z7
9eijKABaW4+D3nLE+eZFKKs965QJiLpviuQQzvUluuXeSUjz9pseCY/eDx0DD6ln
1Jh0uio+z7bCWdxDlnSfoOwH/I2/A1D678zSpi8+SJ49mxa/Y+uIJrdxc6KnVmlP
7/QExVlUlK7Ss5/2BKHoT/mzetXFfbHC59lPUPTQs8sX2U1M3bCPsKgZfWKdYYiM
/zgX/qiZsyooNKwUgBdGk6FRUeuCjp5JxAM55NjLo15eF/9bfj+uaMp0qKcpsvLo
zdnFCMZP5QD4X18HSlaJbubdaVpze1DKM4BqRfGKKdTq6WdDJtVLfL2LLGQWHSOs
32WacH4eq/n/wAV6ih0JJZ73rlfab3Gi6CP2EJkq9SFdR3QFlHTKgewzQNc5OSDv
2CFpPEfpN3wyLILL8+J8iueEJpYkgqAAafBfmjdBy8GhflqJ02DAFwAWnlp3r0nv
QaXN9mL3zLNIbYyzKX6OA98bnhwGEaZ2B/sA25FB4VYSI9fDdjd+KQoLBhkrYADz
f6rmq4yJhrlqDgDZBXa6xNlvepeYNuYPVzstVhpu+MUPzA05PO6LrfJinYJL/KNM
89UgRQ8C8eAMAzif8iWBzTkSCDgYYaybyGmd34EEQtef0WqtnZ6Ydre3jTgxV2ne
nEOUEcTErg0Qgqmeh3koXO6DNga+Oa+KTr3CD+U0tvtRu2rSuyWXeBYsRG9+aPO1
OGLnAAgWda3SBuoRRdP3TzOkdekfDuoGgDvuk7qUcicAyR1z3CG33uMpUrxak6eF
KZXTAWFzPIHnjF1CixQJdRZk7P3jLb1jhgiRiHYBjk7FkM5rgHBjKO8W2QOmcBeR
cVc3E3wH3zoXW8F8vsrXHqXKzPZsLAp9MylVnMgPnzOOMmDyo77SmhT3LNj6eELb
EOXI3/fbCeeZRIWzdzGAOqPDHSSnStaEGtSJ5eq4KyzC31cHACta5tKMEnPlANU3
ed2cf7qBNka2Mq2cSk1d4DV/H7jWzPOvt9X4OKNfBgDFkaWc56W3Y04SKb5n3rhc
KL0nfxjRJh4hXjiNeASx24SK6b2g0wrZtX4hMqPDrtY2A+tyNmHq47mntlsz8Jlh
wpgyFZCNKo4mNDIao7g5r9UE40bsjnlGn4+YG2HIZrRvdpTx4PQeUWD3soqUpaeS
URtWDbs5dK97gQTLhVmV4/LK4wGWfnKpgkwEkSWYfvCd4Axi+Mkn1RgaO54eVwq3
lNVGpurkX+Xpsfgf5EjDXYqW9Sn6TGYJn+kPyfy7Lg1qKO2G/hs0xZUdTXKtL+DV
Mf5CGtRAJ87iF5wtMQaeaYUiWPME/FqPvdIW9zzzw+j4b0knGTCcdOi3LEy8HPxw
aYinh42pUpbGyVQvrC/KGpfgXKcx9Ovd3PbRjyxpcITzHgRuw+C8nxJi4UzYj6Y6
4xL5h2E4vVmNlMDqCoQd8j8HVAdklkIp8+w2oRfgfjOHX2p7p3gzt1d2h3mx9i01
lsT1SnAEkt5t76LYfUi5BryQGRDUnIkgdRWsF5bMm8alMcJ7QZmRjP023Ow3Bult
8se/VDydydSKNxgbeHp0eXnXSdzdEnemz5JGGX4W3vjwpyOctzXnuNpT9DPWUJvD
tn1PCPPmTU07xTwJAApz66KRKRnl7p9nsfQAZx1n/f8VFB703+JFCAFsqp8v8Y8Q
BjzBum1hvhEn53bPs2k0lepZDtmSJ+zwCAHqwSAE8eyOgBIKCMfxGA8V6/ZM4EWn
v/NnASzfwdinDlgx9kGFHTyJhU7S/t6HtnQ4jNVzAO67jq85Kbg46kDNeW8ttB//
UwNC5Vn0L/EooTwsCF9h3oMyXTS1D6WtOnD02z2zSo+TY9DL0HNIc08lEOd+5Hrp
zucWmXvC2pEgba4mCvBCsz6Cmr/kiOrzuhmX8eFSYB5IjihxUKAPLDLi7mosmGq+
+XGeMhsnAU/BEEn9PDTJ2EWJgYi8sE3tWnUbqbeTgHAVHyKpN2fW+HpNOqOVv/LG
YLuS/LsvVwDuu0qOnE7UMrVwof9is2oFJOCxdw2g6m4BBRNbIbMA3hRO/HtlyWEb
uMviu7I/rz3LBBU1sSfGbEPMKzk8GQDUwOUJGdDEvEs3NbLOiPZEN/SZ1noHK6Uo
LfIU2VmA3VhKpa2IRS/XTFrsOD73hk6lnVhRgl1UYhj8qCswoItVvTNt519xJ+kr
CEwlc2rf00EaFsfgDPPWwB6B9C8m2dOw3B+s2SFWIq76v3eNEbV4UnsBhdD7ApuA
L5tkysdrOt1dh+FbqczN8MECdNdlsTt3p9zy9oPBLa1CQM9pSb9tWHCk9hq0E7/F
5vOjSyi7O9IMFHdeZtpToGlEyDdwG93ukHt8l9T/25tA9nKYQI9GwZhezSlxIQOk
AD5Lw56tC22/+roS/xXO/joSZvbDNejpTEoX8lxM0YlXkz5G6qJMJVvAGmiQ9y5I
4RuyFwK1TitcTMWQMivN2vmUwB0pODCEge2M9igHkc3Vf8efK6zS8lnODcwm7bJt
aob7UPcexNp5nPQvu1R8lWyXaiOmAbfH2LYSYImzkbBp/PckWDCvnH2QitvxBduJ
lBkwK6tYQfZ1tnMMnSj5Tl++lqiJ7p0v7aQMrhpfqZ6q3gfNARtuJA6W3oVMBp8O
h/1WbjNy1mxhyHdcclbetjH/r0qgkzGswEhM7qyFkZjALDFIyKWTGb2cMKNI6jXa
KniY7m5f+BTihCzkLKNdSjDG5n6fo3Q/DDLif6ob1fIkBh7odAd3HAXhXoxSaYRb
jxgixIP5Ty0Tt0F7yzlRDRsj1WGQbE9SZy7UTPcsWw4lqQ69ZG43gVk/XGUnUSPH
vF53sNeY5Y80bAs2peMIiv1dm4snRICRrpAbJS2gkCmtJPJbTEcEgi4N9190itjC
W1Uof4jVFmqiZW/AEp7olXLShQsBt+6aqw15yiEvHGHULoiqVt+uhYy9PuwUbejd
/7nQEMsRNSzfDeQo2L5vnxIL2boKcHV5BrOhZOmI7G/EzTcTaOgiP6u5HBGELcII
dA/RGVppkBkchFnffqoj5B3PV6RxJVfbebFuiSz7sOARNqpN6Mx2NeeP2BLpvUz2
f67FIEPnumuCW0HM/8hAb0Azy6zzG11yIRea96a8dNlWw5t9ET15IH5hIQqc0Mgk
pagXocT/4TQCcKaXnV8EUrlpFnsGvizkBs9XL1mlVLLCUn8q0NWI4YFooduv+hCX
KpW5h/lkN1B3HRR49bKVC/hHZju6Xx9+4/zGMWGxf1GCC0ZTxunMTrlq2VBfG8a4
5mV8OUqu5Nmi63c6kMJBDa0aE1hnAHeXaU55f+wm1OEIUXjB9/4OBrjUZF6ezkCm
rcZ3xaS/t7WAltx7sKPTsJBKxR63MWKWQ3CsNc0n09uAfajrgv+yDqgk7D0+KqZY
L577nxicPisXYoVsk0cic+H8OdaqG9deCmzQFbl1PnojaWWsEW0EGp10SOL51ca5
sKVIE2yUayyb+/PuosE0YvGuMrgMavItKXhaScFfOw05tWiqsZekgcUkCf0ZovfO
ukYmowXrTg3PoTwhT8Nc54zuUFXF5J9g17saDlbz8fti4JPLN4aH2RW8jSYON60V
cqMm975APkISm/fP4kdrqEOnd6YeLeAOPMXWClfsuSA4mfI6fHATgzn/ofnKdYIh
Us3OjZBSaFYpQ5E/UfNh0ADf5KUCwA99aiWmzccoskfMyfM5amVTidG1lAJea9/Y
LY9uUTJSOSQncoc/4X2Df6a16+RPOxinLomT/IErzt3WUJQ6Y0PV1LCrjGjZta9E
SmD2OEdzq6JFf8/dJGWKnCuiArOSe+mCBqBG9lsj86YFjf9kI30UsE000tsomQ4J
GGzqdR9qZh3qlNOdN49hyfCkYyDjipzoqx33pATbRsrF6gnnRWy8wO1TeleE7OA2
2TWN9Y653zNtURinlqzQgkYnTYQ/JeQe0KH1N0LJkFR5g2L4InZYSMamHR0hK30n
g9cWL0hZJrGPFS/xBeT3A8/jaINIQ1QI7fjpa6rXgFeYw0nVKFl3iJZbjdzfCI1L
Y2qZHAiXVCFrLNqe/J+UqcqVZT0z66vrAQ5Mf5I4VyxZnV9kNoRkML5855Fr6jot
dSlw1z0wELVqUH3yXxLaPfvJWdl1g8yjfkEeWBMHWK6XDxtW/u/zu+BAV8Ip5l/2
Fm7LgnQRbXZXfJZNK+gR7UTV2tPuiAO7e+i31jBIriOaQ2dlaJbgxe1pZSxR5nbm
hUU9AveCG6ASnZAbSxt4FkKB2yEsZ5hHiaTbvVJ0mFosUNNtY+5Blg9xVvzJX2Xb
P5CrCtOTao4vH9vW7ARteiYcRkz0EunG/uU1iW2/8lrOeUlP2NqiTIj8Cq6j2t1G
ed1nC0yZTDeWzWhEhhlL0HNBEygwYgPJh23J3MNefUH4ZxAn8SC5A89OPYR0BFfC
Ayc+ihKWMnpbvdTomY+U1N4o6Q4FdCNHXe+uDaxMZhqR+jx2YmDEKu+qj1MfNWiv
8k1o1Ql4CY8A5F2VhiHoF+zAZ4+By5mv55ycnzRxTtG7Gvx3NuvlUca/VlVINtQH
PRhA9r66DfzOSC3dH4BD2UX2ss/0VAjZOCgjdjF4+MQ7S0u31tdPJzjRxWYNgRUb
uOXA2KbLucbZAu2B0f70yqUjmbcIZU6r0hAfG3k0wTGpNSZ3ja7KI7/eQNCznJMz
zMB/u0MbVVmkGS0ivO2i3QRf0P4EaUZ2CEM4yE98Zf7md4IFQe9Y/yZhXyNaCgbZ
88R20LB385AIVDMjTYHfpAWKvfe79mxtqXxH0ANeZ3ZC+pTQU1p7kkTqzmdzVhco
jNP8nd5vMhIHUtu3+jTVCd3wVsXEzCj1nbTjLwmmE0YrbU8K+ZsyztKK6DHRIL1C
lZdDQOyy7wzSC3X2jg9q0a0Wfbq5LE0j778cvig7NHeSkgwiHlLYI6hvVmcOAKJ3
a253H3VsFOn3ntPn/869a/2oiUDpTnWqa7LlsUMs4kcul+TKqTy/8qiWi7bHFQ+B
o1KZ6erbcKdjR273IwIvCmNLduf8Y+bevtImQsE0JgghkFBlyiI2kMmLcE9wWJc+
ndaUipbgkRGcNIV0d3zun98oPsTWl/fxQEDMswopQcNIo4y08uLKgHf3Bgs4ZPEQ
b63Abs5acBh4vIqG5iMAKjAdJSPH6raZ+Z6lNpDEowe20IoEKvxouXSg42lutUgM
oRxSMaMXFyeBtdBqCw708WamaPrL9nNUmQ2pE3sFwOTsMoJfqhi0WdU23CgNX79g
I9Z6wSt7gnMV392Hgeg3MQ9NNigCrU7H9j34zWcNOUu3sVdrfBB1IEVq/HXFFkgS
ZFOYRZkvsx8j0PkQQmve1VkzERH63PJqUDCKfuaEWoyOY7umtQ+eT+xUIxh/Ejpf
zccmOV3cOxFo43D1cc9qPoxAI85RXeENNeKUUAWpTKviIR0mNh2D5jDC34kIjO2H
XHUW1xkmNFkBy1HP4phCZxh4WYIjwdtAeCbImmcX+Qgjbl4DwxYgDPFKwHWM3aJY
36kb99VKVYADSoNGFo1+pmqnQJ9kIKv8nY6PQMQh3h0AgnCkJ2lRIn2oSwSvwZ+y
Mh9FAsH0xK9ZckYeJP0aRiI7rLQypHyituI8yz3ZnV6JFSxiaxjL+t3qgPrDp+3o
XDNO3xaMs4AvV6oM7RLcsw6bRgs/HgLH/vbAkqy43JgcktpatE4lo6Cr+xmYMqF7
Hy9V+AOVxUcjhVhD9bQDFXjgm65pUtS3KsjQF+5GpQc36gJS845l0SPJCdwMPaX6
cYIpjl969vAFN+u5rtiYQtOpK7s2Qv9bIid9+Y+Bx57nqlhWnzlLtuzlUxVMyq4u
KQj5uP/avSRLqahzo/mV3uw1RMCw2Nf6HlV4nQc04rDefgglcnRNCL9fo02pz98n
HunEjeJkOULRZ46enhgvHEJdEN0zw4PhxbXjOz/VZ4k/TZLJjRizl0I3a3J+IFLj
7G9epV4KBw517jzDYsCku8ATCgY9nad0WtMGWcC/TSYtKmSCnlGVj7zvI5aEv4x4
9z2XE9lkqJCkmjfy3DKgdOFA15VDkg5ffPxQ+W9OTg/ExOmyZd5e58YY/22rb/I6
nKizmO03cnqoVojDit0Vji8s8ctL3bdEwe3VaqJY4WkyDOGs85PUfltFQsq7SoQM
ML++VB5QtYLWfdodPA6Cx1u5N2sDdD91GJ64xXTdrNXtAdtq1tVy0whgujM2cl5W
Yb5eTYlM4aoVGzDFdIPEnM6CK4Q8Tb/uy6Z3sn4dWBbjSDAgVgkVv29w1gx5C3XA
6d3gTLLSIPeLzQHLtKK+QZyLOATPXoCilZhGDvxov5gYgVFSvBxG17a/7amwTQcz
cwYOLljNngnajM/oRvLKEHr4z8GUQ/+ipqA9pf7is1d15+Y5R9a3TcMX0zyQ1Lav
yeya9T5T/JBA8AvwHyX3poo8Guu5qYoSatAg2+xG5ZtslE/IiREDxoaElq6hZGtm
3fK6ggfc0AjJU/kzOOdcASgcCKLqT1HiJEOSwEKocFO3s7BzGPtR9QDVdhMHk3U5
2ly20grJV9+y0ACNtj9ZGZy3LHstncW9H/GRvRvztvEso+TuAxZgnrSFJmQhDnAh
+nJPRkcmLnwFwv62YU5yQ/H/QsK2VuM8gmT+K+FytPFRJzIR5ctnjKaAMInPi4sV
fnmTP+rsqr77efhoCGphY0kAEb+4McvBlEdtSvg7YcqOiw4BMuf2dTN3FvwU44QK
rGSS0QZ7QIwU57f6H8ZGAB1ep8s8v0GnVyxKgwkPZDFpW5ngE9uECRIXCE4ti/SH
EAYWIhOaR1mfI6P41zr0v2JG+fsEDp09V62XyDcoEPXx8k6oJCKrt78kBvCsQA10
9xENYuP7HkKdfOkRS1IsUBI7JkL/hhnob8o7G+sg1HvUIIu1zv4b+c2RhE+0XJ6D
Z0P10wZoXDXFqFDaulJaNR06W4J4226aX1ypn1CaTBd3MF8K9Qdd5klFZ7ArA2sB
B3pVF3U8FWoBZK6CC4RV289rLjFE8eyd5VyP0Ph9KiDKm/VtxTAoKo0NYZcYv2ep
0OArfSquGkHoVFP1GsnnV6TwC40jNEtIjsZ06udHmUMGV9CrurSSasH1egUUx0nR
f/ElNoMjLr3MEgFu3LaekN+LM6cmyixNeItf7KZ1Jj9LcDvOPFpS502imurwJOTl
oeIwKJrYSphvz634uZlzlTS0XlYMiH0L8g8LE93BLSHTjk3WFnVuD9v/VH+i7Bi7
noFtmRGV32V+3zMlA5vCVwWw6VHBLlM8MvhZAiXghxZnSfBhGfySTFSSjEMKlx94
SPtk5DUmGuG3QhOj7CQBtL58D5CUM/HSx8mqoUNoNI7puvdTTbmv3M34SokolWpl
D3pQiPKXoUyjLlTCy/bjfelIfo5pdsmKBTnDkgNhJrGovjx4JFqh8R6Erf65oFLJ
YTULc/rPG6P+0RnYXI7HTlj+O6pGMkN6LHl3wfsy2P/KZ25Bi3HvYXlB+Rbcl+jY
kPxCek730yw63OUAYTa9wH4K4YJLBEvzp6VzpVJwK8TbSTWGiHV50n0KmXyO0tWH
GQNKOLNIqeuQk0hK0Y5MxssuRDJIbHOeEus11oYexyT4bz1tmyDqCPDLyC92oV9y
ZnhgaSaSAZYDsKk0KppaFcJyLBGH4O1jd8NrqtQVugA/ZqcOkLluyGtRzugcYwKw
wE1XZUh6QbKg49ZE1x8NSDs6MXVYXw1KrPM0tWG5r8105P70bpbi0zie1WPKpxN9
DtjhTD+HtFKMGtw+5+IUq3SrHAggt3BS/VJiJ8Q0XbDW1WPOIGHu2NB96KyWrRi2
+e0ZL+aFPwaEsSsZnLu09J+07N6DcQeg/Pi3U/dWE90FwS36Y8dJk34ZsEv1d/Im
outDPrPjvumg46eJ5mzp8TGnNO51FbRbD/VEAxNQwYdBzz807O65jZZx9kGRIR5f
OeDqO1kIC3yYnTaW9d/WEyTmYNcHJzIAtwU4hwCVcSKow9/dMH13IqFxadlRf1aT
T580VRgmp66/RIBbYVGlhi3JGgx34Cn4s0KAD2I8DI08QJn4qwZykA4BXFP36ZjF
Obh6sVfg47gyjjlM2nwnAgxJbxmdGJ6uDOAG42ogWbOvFbZB9dnTC6xtqlUND0Ql
4vLdabPyRaEyhVsnFyPeMxpXe83Wi0nHkdM9/8rtuHvb5ViWLnn0ntjMB25OjxPT
m0/KujDNSyW4qcq1/nkxEgVYQNpgMCMf5PuewTUGzoNTnfBWAVG7Xh/y7swRc+Xi
O0wSLBeduSCn9YHhSG3LqTtizl672GVzEfCPbGhlIKZF2fYEwLmCyUEwm1vpjO5H
VZZZgLTkS50sHe/dQU89zST/rXaIedR9sK+yDtsPOfdd+vZO7txHJ1dKoVr5HvPs
9NCn6yu1BvI/CcQYw/5TVjjxIljgW3seOhiWDGf3QuEo7Yi+coow+Bn8+PNpcEJP
YPyOF2oI1LqSo9y3bUtMtwZKUA3zjpP3sXZnXyIhF77qL+BBuDPyObth3/Eg/t4U
pRaKT0qEEZabQth+822YiuQQ231YQMZwLM/Ya+qB8x6VQN/OaNCyaQyO4Z5BUdK5
EXTwlYzJ9+SQosFVpeVTNSFPGeYYvx7SJXbO8iYTA3b5/QNluuZU5sBgz+F1fy/4
iry86pRZjCi+EMKVFDS4keUwHmh5D2VBww2MmTi9bzAOiEX0lmpMSvkUwxl5ax5j
uYGK0m0Gn9cml7RE7iv5gXLiJH6f7PonBsnf6pG94n9n8UPcnaiEemvya8D2CrcP
8n9M7CULUfd2/MMJRO+AsJEapzb9VB8CJvKavAZ0tPwQgOF7/bJkWKEH+IY1OK7h
CAeAUXBNuK+ve1kWd2hh23loXaoq+/TtRPnHPxDLvRf0423qZkQLITjfbtp/k/Gh
vsulD75GhnTvlhJ+EavzY30WSKV+EN5h6MkRlwxhSBXM2iNJUx5PwY7dIpf4/m6C
fiwNOXHNqrEmGRScr5XPGQDTAByX9EbNiCSZRA21yhigLDssBIBsOirU32D/6WXH
xDPB8EQlMeslzG4B+BRlQVQRBEwjZs8oGOUS8clAM1fDwToU60fIc69R+WsEqxNS
dce8LlMoDTI3Go22gbTCbXFN5jNUR9dW+ugpfebSWWO34mHGHgtfsu6rw0osSVyD
T8ij38eg8cT6/lu8/b7wPiosh5hf0qTDA2HHS67NkRjvLQxzVZ4iZIjc2iDY/FHF
+XSKDDOT8bAPwrfxuIH2UP4+4sFJHaI9PG17CtOdrKZRwDoNYvA1T3zAXoODku9s
SyjYi/4yOXztK8aaRdiRiqaVBzlwAqHevCF6VjP8xfQtSH4HutHYLn2DSM8F7h3L
zex/Qv4e5ORrIOVGT50l/MZtwakDNZTEE6ZA3GRFHBp4HSLJs95odilIL5Vx8bmG
A/j0LtdkNl1OaNdKV+W51D78UuhN52w1qLWbF57gdIWnm48PL/FL3ma4ZjL77XCb
Eb70M8HR9CV13gNz/CfrUX4uIizi/o7Ohf4lX0e23YErcxKcz5bfOYjrCf9/e7Uq
0lMxm5vrRYSWpxpUF6pV6bN++9XlsP/IWNTcik7ZBqmTYV8RMBl9suXpJFgzPkb3
MS776P9yoGtItoe2yxenhHyzlKEeVPVUUEmbqLzNjOaF1gqM1HmGG0n79tcFQ7Ls
NUmwTRCBQ/txUDgvs9JlBMlp4SpQsXjCH0h+gEVXkmKp5VCB52pcjD/OMTlNbwya
He1mpv0NHuaUGMecIbPlEUAqZKNQvoE3yPvKXT0bljw3dySvjO/vljrraTwbeRTD
e0RFiJWdaqVldK1jhLMdHHdHWXIsvF3tPcarbsvNhR50gFnRrH2PzRsfgk1q8BfF
5EvbE1T//q1H60z/FceL4WC74+p+QhgBsAgkMqx2+tEmOnJokTBwBpXC4AEP7fK+
NVmwe9e9cS5CsKg+t5aooDIMJalWZCkytSGHT3VfXgZ7pYvzFgzyU6xhHxhnIvT4
jU0zhzLfbRh9ddS6uTeSU2qJsO2etlMV69sPoB0jXxhjkcc6eh/oHC+iYadNTIzi
ttZONlq3Me7egimRfsLvbJuNkjRaiJ+0qyRWPBdoFLX0ck6+IAfghsAkrL5OvonZ
2QVrqdtr/HdwuI44zxhCIpvHf++JBKWXSWl/wTxUhTym4O/oSjbHMFYLR/vNwbVu
XMnti6HX+dPPDZG4WXu6rPDdC/Vrd+flzSMBZatUlsfzctxLmXz/5a3PBCmc0JNs
5wUM2sCQCzSIOOw/fXiC0XGkVtYbVEvIYemIUdC+iDzCs2ukd3oYle1bQHnEd9PO
y3ItEQRUUZ8YuDWxslRy00wwrXMcaieEhODa/tX0l8lnh5MAccRKyN0m9MLYeMk4
rxn9nbsjZNjjxS37WA5jCDCT6AVld7shqRCAZ8pvJkAlHeS2myBLCPH/Eh4lSWpK
AyDxvTDhqBukYlv4yibdme4sjHN7jp+z8y0/ktHf6BbHWAkuO8oOhqSGszck+4lu
4mBBrBeiTQUyP+CtOQfd00AC0gS3aP32xlaG/eqGLsaR5s47eAH1g/ECgBjwKdKl
pqo685AlFGPTgTkIpDugwUpr3WAzr5WdC6eMG5b4yCUXrqL7iAlvO7t1QC4JGl+u
JLLhWFmHYo94wh5Et8SESfpAhOavxJow+1HQfGVBYwzHNpzQHjb/SqepErKamnem
e/X0MpsB666CibVDWKdzKCBZFJwLzaQsHcLyf4OPlYam/wLfZS3iG3O+FKUkYUaD
z00ui5zJnjHvvVZRw0jzqk5Fz5nPyfp8LEGlIJ6CSobItZY4Rq17GHRVSe9hHXUX
+pvpWFMmDh5hRFo7q25Ib/eZJQ/J1eDbQ4j6OCJlpqd3NZ0TG9vb/hT0l9d5qdIe
lECqRHhb+tatrfkw/r909oVd/6skvgf46rlUwthbFIrd2VC+Hb/7CvrTBi5frLXO
XSBWPZKvDKScFFVLFBxWZbz9HMYmA5qhd/vTfA3X2qkKZdtYBDHmBZ2F/c+PqMAl
qs3U7vAapkz0Wzh2fX3sV1uLIfEkJQXY9RtOWJ+cUXOg+4KL165E0ssDYp8cRups
BMHZZ5F5sK6LpIfP8f9/9OtnFKrIQ+6AsRwsB7XhCoonUFj+R2GboBitPwgvU4NN
ABAJKPULt8brkhjlkX8eZ0zCwQGM45/04Yoqv2OliVrHvWDJGjOIJdCAajrkRYKx
LEEnvowA8mP7UX8YiUDAiXE9+oBsEt0+6E9aW0FO2dtjCsmEp4W9ftXfOdzVZ5w+
Wvi+sjoQYYh3Wtelal4acR+fdT1iQ7aGtHpvEWm+cyYo5RXOURDtE4ga9hVcGZNr
S/DdTNuGV+q1PmdzdcBTLNFiHC5WA8nP3EJ1EladFiJs6gUk0rH9cmBCh+hVnkgm
PLb9RraUsbi7lnbfIhUyNL1VKj+BsGOJzuEAXMOnQK+DwJIPAcaWMcRERVumKCrH
J9Lty+bJnOEORb/9yCVfAYu9xo0yOuPgsEiEUVbg/dCP38yp3o0kukFYtB+5GrQN
EkSEGcpoaEyiz7dDmtlpPvkzYavSQNf1WWm/nFsnoTHwQ1SBKP+jopnDdi0iW//l
JvaUTQtG6icyZb1aqGc5hYc1ElX9NV4Cg/tTjlz0jMXeDwfZo96tEOfu0dHmM5l+
dqP+znKJo6UxFJmeqKeE+7EMLocf3Qy8essUPlyYngDV6PTLMDblAHJLzcrZzBfB
9q2d4ULY5DPQbykZVdJJedIj43Iv4BlGxOAZ3Li1TVxlZfpl5LY26nuU770H9OfH
75SEYYNF3AhGE6CattLUPHi/EjTcCIC7RP/xY1hFB04hdazNNkYU/cPHNqHsTxpi
pHBMPAAVHz2VaNS6Y2UNI4XmiNNmYGQjM/P+cqR1/yhk0lD3NbWqUzpSJR1ByvPK
1S78NS+4nZxeHk7QSkPPN1Qycxrh39Bk1k01FpIek8aqkHDWjMvgj4OXpy1saU7Q
76Abs5ivKL9sKQZBmv0pKGELRKDv2ort4m0fkbT6hL+nOPyLG6tIk4Fp2vOw1knb
NrcuyY42XfLpBPTpOZBBHDdf7CwSlmLZkjfqivX68DF5fZAaSKjETk4tlMtylSiN
ykQwgeyMgptNktrzY09AeUE79ZwZupf1Nn0AFhrEdr1a2KamzFJxdHBpfdzJENqw
k6Mv37RcFRwbnOX1WTU/Pe035FXZ4APcTxJlKUTZewV9ZSvCLF5cH01JwhvOaAOy
BJpRe1U2Kpm17RrsxJeVdCKCC4BFz5lHuLcH1N2KdHnhc7u1ubgpHNAVrIpPyWcN
JXG9p7CQ75wmYGP+g1OG8ejS2nkIQt//+OTzY44xAbFYZ0yWTdQ2u7lXnrqmbz6m
vDN/XC3bZ90Rz7CftAOAAOHg6OYtVJ7hf0Drr7/8SBx5EHWBLPOv0sFp1ZTtRGLg
Js6bL/lr7OwdUnTI02CYsu0BDCSmc4AcX2qhVlh63nHmzinbg1r2dZJc+LNC/Kil
i3MlVcPVbgkp6My6p1GJKH5OQyYBi1FLgLg89cXgOt7Mlo5M66Or8ojhyIoUch9U
OK7hhEjimYBQPLJn9PATam/7J6O93emaCQ2yrgTilwtwzv3S1PVl8vjGmTJM3rjo
7EfTfpMuyfNwN9FKysXHRRrU7h3XsjsxwsyB/8cmYnVzYRYbXACMqHCybuuk5mxt
w4Vmo0M3uTRGls5BKz0DmIhuWBfNZYTaB46mtTGBkLtFmoWfjV+DPK8b9LdMqZCA
scshRQtsze8RpR3QwfGiew7wYwZhXCW4vmp5rAx+My4v3q1D8WKBQLtF/bxtxu1L
uj8Cn9JGqKYjzANggarPK8Wa0hXy1RafzC94CdtB88nPTNTc9f1zWgkVD3kMMd81
LC30Re9tFQvG6cB7AkrzmIUKRu8JvYeM/v4oTJWW9BfdfpGzWPQ6WwCVa00G5MYD
4/ooJk28/YebSLZ3BnsO/Xv3Dzc8d3hm5xSnI/k3h/BMN0MuBliLLckbtfy27cL4
Wk6jYskWHBULp1D6lnVTEoD2Sba8wcTSh4oNy1XIe0xyYIF4oBVB3TKq7l3Zu3mJ
rZITung/JanRFGjEUw9MNrb+zozKOa1aZr03VoWaAkQ3Sm3wFd8cgHdY/qWgKLx3
gcEjXUGzyRdznWqLPDTCSUXnUF0n2Ic/BDCIDeITnm5AcXb5jL5CKnzp6Nkw7Gdz
TorAkOO6tCL0ofIDBbyad4PD9GhQ+7XB1x7dVuMZD/zWK8WZD26F8tFTyIXMorTT
JxZwabjf4JJEiz8HtC59el3f9t2pq2fhA3R5S7S1QkmxS5Y8ltR2YMV1zklZb83C
2fSJJBLkfT+OjkPgibOcGxdMPCa9C9Ig+zUdJ7KI5c/7ghN9XnVxueI/lzshji6v
dont5W/ZOs2CnhsT2tyXFEwgQBBUWdLr3lb/Rhp5Yl5TsKFx22Wp+v1cNo0syBAy
h4vRy/prgUc0Z8meFyI9Jvvv8yXKOaCpuNDKxYVp76HC2bkqS4Q4dP9pWoQiDUrz
2j0Qcp7yu3QSvN78XlVM0Xpc8j2iRyfUJP8LazEsc9WCBpjNtG87C1RkyK2LvNNM
vclLpPcD9hTnF1biZz/pIZONR1UaIejYcXBrJ1QFxKLqLWYyMujAPYMmlDn7fGmo
Ui1PLNrn7hAux6CxTXukLjKLxq8P2cMGG8IQlD46HqwKfXT/CBDFdBGiZUyjaQgW
1vUeD5eoKkdxzjkD88Hg9ikDvtEhsy0d0g4Mes8EAd1PZZecXD6u8T+sWv4q+9H5
2G9ieKR8sEgwgQZVaqZEz4KLdHuLjEFriJGLt/xUVEY90uQdK810CHRjZxJczCwA
/h0e1Hq356vipwxU7ig10x+xvbesw/+Riuge/Kbhcx1J/3Mtfkx9p+snjsP7BLm/
Jjd42sJ486efrTOiP2NF8VraBRe37JbF5PEpukF7vCELz0wuKQwpDA8EQM8HxVcf
zNr7OxpkWqa+AkTe88Y4nMoj64WbBpYRrTvD3Ht+Z9ez7L69M/HwdJH6P0DfcS+h
x3dd48ovKlVajoYShaPV7a13vsyciqJ6Qq2nqlkB1M2hYKUcYjVkIWM3vc7iF0EZ
ATCOIDxhijitv+efsYIL4ANpF/Bxj0GodCoUxDfdJ5cKFjxFdvO1UvCy5ZW92Zsx
uEiepNCmQOstBpuEbmOkFCxgBCnfzz4QMHgPJSPHAu7C3cEp1jymu9Gqiym/1OAn
zx35hefFszh6nTrQHakxK1WtPQBYQHxRZ04z2ExYhC8ui04W0PShbXxvhJyRkgCT
7WS/Svy/+Ec/lKE28N992iXXLXTYeKwrrfISn/VSlhgWkH0qo2okgWkg1S+JOaRW
FB5SjwFw1WJrGXqTVVENvFlyloaw3mOyyYSzHo6qRVnIC47V0bW1oBp1/7ZqaZ0n
MzXrQuCdG6R3nwWEBnOtiqO09yBCZ/TZMK8++fw9maNYWYupIvnoO+l2CEvMxbhg
y6tmMNtof2T/XZImjWiLEP+iIyT+HezzubVdHtnX09VyJX5dp6OcANfmOVIBF6rY
1hS0+KHZpuqhP4Bxvs96sFiN94rC/sMWOxYzr2Yy6IYgBUCVPhV89eGPbXEzkgrt
mB8ZUI5nDvjrR67/pPIGXf/5YYjIAN0NR2cTI0j61zatjcle6iuJkJPfUCNVQ1js
0/LR7URAZhJ4ubdpd2+2tlT4ijFIItcGWzAfp9qd7mK+AlYtNhXqNw4DPCTtbIqb
bqh7GjlBa/MQTacixf+YTFTeXiK4qK7t9Ao64qmiur99hUc3rljkah5Og1RwxdVw
0sCI4XU7MSAdj3NGKJG+b0mSL6tf6wX+u5ku/dshqbJw9pTq4XyTk1ZiVXLb0nQB
vMUDYnoV3pc4cP9VV5ZI92GpRhiDuu9Veh3LF/ZokecKGN7PZ+kg1QqeoI8vsTol
Wo4ZqvRGdKtI1YsI4SerJMY5NJqu3JK2QPTkejknL+Q/GsZmmNaq45yKyMKSKBz2
0cerygGQeATxX3lCdO3fPiBMPSl4lyA5Ju0aM33fCZxtSXWomeZXz6JOtVPdz1Nl
NSDDh6UoLFB+aEEYkfqwsyMdCxwBMeGPbjtyu53YHAndqehWlidLR1OcgE0dc3Hs
Xxipv0JzcJSlA4oReiCb/WHREQXUdiucqQ3ueVaKdVbBVQpC8vydjbA/lqvSdl3a
gtaV1uf3kXZ8NoCsxpKfxsf86pWe49npxxtrUb4zq7g9iEvRtfYfATqfwNUkCyfX
gej4ngezMmP9ocEpTlE3Q3yAvRZjqrWBksQQX9+qn9KgQDlyjcwm+JTxNUwStZuI
9BwKuzl5zRXLhsN/B5qqqL3gb41Dm6+Lq9j780fdA7xUuFplmapcZcCSglXG+4B4
ME9uvk/l4uMzbdHYRxitTlvWr4dvpkRyC0d/i0jc2Gw8/vxwEApFkQLwGtcS5ren
j7Q9vj125Ygk1SltqSybh4Bzm4oSLThDg1FobXabY2kcAO22ry+5oNKIRZflWMZA
moY4OylUoYWDOi88CFnpwcnGOZAr8MlYAaadnWX7ogMk5xmXpPy/gpElK/OYMwCD
/nEndYg8cOQ8kIN4IY/E7sMnu6VI+mIJksVqW1JoJPqkfNdzOuqPLH7Pp6U4GdpS
Z3By+tT7cyBE86AhzCCWdahsYuqnsisBiEbmU3fjp3v7HLpa28iPB3IV4iD10p9d
3kEyCIJSeFwQ63ScPGm251oIhY3YdwyLFtERIEAhfosFOuBU5U4HNFdVLezVn49u
n37W0pOWC7hw3jWzgIVHaSLKxD+mBvHPTVrn2EyxdmJl94E7nqLobmjZYXGWhsVJ
ZmEoKUJf3E4L5nOAzHHb2hIrwKcPrYOJGm7zYvcreIXXvOfcM8z/amsuXsTMBjhC
Oh+VBa47ZVw4wemNjS5iCYYv2ScJLIMF2oRYCfkNt09pzCxgoI26lcBplM0F1IjI
+12og2P6+RxpUAGU3l3IqNfUoiLFgOSeDzdbpVGrc9IXzK38KBZOWqD+ui34/Sfw
aiRK7OBEQ2NXKQET8vMgFmzDOq2fIaVRsgotsP+qGxa/M5PpxILrdGLFFoAqQJrs
dPcpCqqHlzPXzM0zqVROWtknBS6M3URmxlMbTIwrJjUVLoeR2tatCSkjzjf1cTn8
BbO1x/TRTajwMBG/cR8XdSJ2ssAUTg6agl6xziUk091ogVePpxjBAXo5/amrU0Nm
SCFbowZyegQiTFKir6UjVx7TgEUqO65O3D5RJWS9kOPJ1AwFRGiVlrcXurgGpyjR
FAw0P43zO7p9zChZcbEc70qaMbDdqBegogHdbmHLtiuPRCP4EvjzUKEXtrlHJK7v
idTrx2lOMETPLpr9k76tmyb+QLnygvz9GykP53pHKbX78gZ1brsj3UI7UQXZfq+7
5wTdJZa8n1HF80A7zRFbh7lUTfWYGKV8XP/iF3+EBaGJ8e4ZAA0/jTiaZUGEk05B
vA2zU9vmzqizpPz5ubnaJXkpzBjoPHeadZo4cEtr7+A6QI6mBb/Kohk2f4E0AvuL
iLXZXd6oqsIOlIYqvGbxn+fUswHiBdeF+99PdyDDjX6mKi0Tq98ZdXURBEonnVUy
4tNE5QUvmm+GImFiC5EkecUAua17yqLY0VnTQXKJrZOlK8iW1HGltdHSZrqzm6TR
dYmR1aHTHDoUjqpEobGCkKtVWCD1luvzc7K1waxAHwrGB7Irfd4kIAIzOJT6N4yW
fVX60wkm2oEHz+ZofMiC/yqVwU5r1Mgf3DqmDfF3HukF0dEK+yJI/zEkgoauBWfa
vtG5LJbb5O8B6Olu0LX3jyyLb8fi+Ah97illF6g058hiC5rTIluoq6+RlByIxb0A
9RRJCUUPIwBIpHPj9XUj3FDnTeQexjk3eDKU8UJ6h6jMRgmVemejxf/tnm/4Hylk
nQOkB3vn1YDLbYfz7zIXQ6B3qIoTVAifvA1QUfayJDnEB2WZd0lx4rLZTUlJXlOi
BtlJdR55PjwlZZasCJ6ifNMIfSUO0wzUBJUMOfXnwEwXVvy4uZ6dHgfKYsXF0wpG
l9wfaERu70kSQMTtI3udqUyy+m8+lOGxBu0pj1rqc2Vma0WTxZ0id8NIJAO+05my
jCSKo3lwHDSspPkiONUhOAi/KDSdIjKNtwlYAk8dk9s5n0WrZ7Cws/IuKvknNCKd
SuKRlym88xpn5cXzBjoq1mVZTYCp7MzbBYGUi8LHTjpv70KMybHuC34JLrf71za0
9vqEZb+m4/Gy96kS24rjhM0zTTgm17XyNRdfpuT8k4v3Pi2ye2cMp+aOd9lZ5Ozp
xzxr6zxcQypHWmVHKcFAPgrtsGN+XZLXzdyQTdehd7U3hCQAxLF1K80M4GqvtSRr
s3k5zO5LV11zr9J1QyjfGQnOgNvNDBOAunX1MPcumQj5aB5koPaoKrsdU8kGwdYs
vQ5RYjrF91EERGdS4SeEh8Hnszb590MPjRNjB+GsX3OwN9WURXBOUPpKyyfM5Mf8
VcoOYJOBRuPGQQe+tbOhCJ0OjMq5dASsnaUTAWHvpp7IEXEHIFLEXmcxUpeEN1o1
10CnbxoWIaSGo1zzSna7h001YCDSNMhVPwcQx/7G6zayL9hP0TmI/jEPVgttxaWY
BKLEMTTpT+cvnokdmYE1fb8ySbYsHmj9KFLo+CrYUHYmNHxiQDUwpFikA1BenymS
pQNoYXq+/Y3PYkyr55CSud5/ZE2SzHWM+odkdjRtPj46n6pOuq6478OIhw1AaIUQ
VP5yenrUkptDcrcIxQYUPQDYnIHH4dxIi03sp6PV1B01dpkD3nUZOXvLyHdgThFR
AVSx5EKK6cP7ddU5CEtiRneQNJa2x8ewWpssn5nLLVderJy6ZmMjHEiff6z5dEYc
kRPCVvdfP6amEiJ7geit+fkezFqCwg/AsjedCMe8Q+iW5rUewYGsn51sRFMMsli4
G7NKGCjAbbL/oTJS1E/MZgVEvfrKGEr0S4nzujOeWmcXggKbMXuWMdYDfpCpPenv
uwfOQ7Ga0VSbiDvDQv5pzNeqC7086oeDNK8RVqTInREYwxwFx0aJoWiuJDka7hh8
4jjWtQ6LDimQa5Ov1qfFNYbQm88oQxR7yFKvcpYVG6A2GpwtUfjBt/V/G2vgPTyV
tfL4+DbFwrJSmMpKvenNtbBe7MI2q5PnSAcFbgUaQ8sCTTyxmCKUqhXdPtsHi02w
afB+JzFV/R6EAOEerpr6+ITDKwMeh/2Yo7nBap3pqXp0tGB9A1KnOSgRRohZYOG/
lc66n775/JzdIT4ymDOU/FNui4sQ4e8jLQteYm3VSgtfBIbRFgMazTf4lIlfsFy1
1zZns+F5VUH3MOfQ8UqOFBi/nVINiF9EONn0gT9vPsTjnSQqEhPabf1r0OItq1cL
JIhttHFgs7siqYNLWjUy0DwXcg0Co1gtxQhlDsgxDj3tujsIr4AB4vWdUptHdOWI
T7hGBTdpk8+ynX1cYPah+3D7texp4OwzvPKWibuKZehkr+dGuhcCukEKTqE5j5hx
FTHJ1e4gO1MdgHQNg5bM1cSqDOmH9Z7zli2UAKtvyNxWomJYyMKHbXmtJjX+89pf
mhcuwHlMhWatXGdT6xv0IC0LK7YRlvQzOaRQ/ckH39DXof3emwAMgroDFhmyeH6l
oN2wXRhTwspQlqBHoU2XuOIZv0CR00RuTcXlFy17Eb9xzd0cbTSAo3ESCs74g6bU
pOKOqti6Anh4q++Y7EG2Pd4X9yU2WrjdbtUkElIY9E/HFkuck4hgukoPAJwhXJ5f
l1QblpYexZDPGYk48bzznqUmPeMEJ6mdmIOzS1rOLqUBwevkmOkQdQgYGKrG6Tgi
LEsQ3kwmXuFdlHzwpbP5uYisdByLOtnl58jjmVPxTF+uYd5PxWCL9hfLMi5TAohy
7OIiesW1Hx1Vm9BAn8hkRRhochIQKj+D+zqVLWoMGt2itH6x99nsyzSmRHOKriXo
3cK4YW5whenSMohqtG8MfV2mqqANLn6M/Ql7jSaJMIm7oScozwV1/jau6aQfiYVb
we2CSpI6B8ASBTwLaz7t8+96PzOkuirGCHYkkffTzwiA3rnz5IwESuCRqxAKwlVg
oJRKlEUnd3zKz0v1TMTl4iyGKQHQIMPRGmUtN3S+uAJhUEKm2Y9/eGApq6d6y5YZ
g3QrJhotIuXcOzjiEweQwEBOHHd/QHJs2zdrQHP0cEn61vB9eanx/g7I6GQXU1Yq
LkKc1aCe7PJqHEm2E0OAipf2BfDLCoSRn8ZK4caPAerMiI1B7bo6TQuFQIElLRhG
TjClqbEmAoORAKd2tXz4WJrjIQYvu2O0ud3Kn80n1cP89BTYEw38vtQs8rqTD8Cs
ECdQuPWcKBwCeKKMO5df0X//vgNyjaMp6fVQ/EBiUtgkxizHe3J/yrjYX6ffwOe7
0TCgflDt8RyilT1zJklE7wc5mkZXeSyhA1gxUV0AFnkzYuo3mI1Qa/bEwUClpHUE
tAETuenVrfEErY/2PIXnBei+76FUPM7znZINl4aI/vVtjbTeELm1T9ZDkgePQJi3
1eFOJwZbxO0ik5A7ExLgLxARjP2ZUHjAcPugqSx8oaN05vc2s/I1bs6OsSEjkahl
7FNMUE7ONY3JsPwXZz7T4Q5WD1nv74cY6T6qNw7rFgirHpiRv+QJ+oTW5Mln0v56
kCh1ct8Db9PUwfF7+Df7qsDgVrC55yiY3pgWTzNC+Lyxqo3fX1oYWZ74rQOFY3Uf
BC4EJtYp7nm2HszgK2YI7IfIGiuckhVoWOaZ+Y9cMQEOBUq8u278T1Luln3ABhH9
JKIS2kFVToHtMzD4zadwwnQFzCqoN1lv+CWlXog1fFw2qe6fsY5eUTb5174KjgYo
7yIGgGO40jg1Yst9mTONaUrTiO4YhcdkzWn2x4I0oXrx9QuQoYbjppVAZZifzGUJ
djOcrrVqsoaBI8ZmQbpSzkeKnQDUlT3SbUbAWIiAX1NF9cD5kLfeFv7ELQvxSf4O
x1foA50WNKFWL+1nhZ5KgkjDIzxVT0V/AlLsOn0Q5a7h7EmtCyVKtrSojwOqq91u
ypHRHeJsTinwE/zgI4f4HFl6d/C6jizf81mny4aEMIZFhO28DbVlXz8Lxp+5KNrX
V1sqh0OCcewp4UvhgN4lK9LDSTAMJaCpcUYOWlpe5OzN7T+/Rp9OFnv30kIlvK0X
DiG1txPv/yk+/zphCeR3Cf7FMImCWgWK1C3xuXyIjUU6HpikUYrVVmIH3drt9j1a
nmaGiuAlxE78ik5HzKN4H2AHuya0af/6o+Eh4YxbstwrFInxbjp636negajBDcKW
fkOuVrs+TkXvSxGMkY9lwwcOM8V+J37wstKSMaWsc4sg6OaVFJuSCf0yhYBlOrGd
Ch90rRwUuqSG5LVKGofGFhgo8i5qNGpPgpdWVxOFIro2aBztYQvCq1TJQCkbysPV
JBRMhBKaZrf6Zd03fSZvdX8b5uUm5LpyVHpgxogx/tlU4qjrGk1ly7HqcqwUGhnX
nRZ9icQYO+GeRpuLB9aEa5oQfpn00TXUMO9+uU9gZA90dpxUHCX5brVilIa8bRlS
I7J4hAKNfCdKFCAoh0H84DzvFwnUz9O8ge6ZCUifqNKA3yIlZvHjeogO3lwM86Mn
7SzZrOtfvT94TS/4cc/QRj88sYH6/NpKSE++uV0s69YieVnLThruQ8IMXailvbNz
eDBOFAbWpGbvGGwlxsyYGNdlPefgwWjdj6bSleyU/v74SuouO10u5ok0rQQQVExD
EevMU19BZjUnX1ppp5VFfnL4lcrthbwncKybjRaDe9y0orv04NyopG72b4QSeooP
Xc1ChBwasUCd/YcyND6rThpQdcd6mCqdXlaeBtw1m2YGWcorQQR9reE1PaYrcr2U
BnvEoGd7Fb+Ptdl2ScTtwzqLEh9lSFcZW7whKeFWfJF54t/cYJR19vGhL+0WzaS1
6SLHSw/JQLiE09f/SxeqY3MtV7tPQSk8vgOaoJmrmU8ob2M+sw4NapwZydGDz40o
1OmrfxCtLH/pjIkDddBwVra1o0we8rbDhWDzIhe7umLMle8bAH++zKtSJJxEZq+u
QEOKoDkzgtULEuaGOjdqqvFeSdVqsOupXoAeQgdniG+w7+RgkQvKjchd9bwxQeE3
9j72eFgKQ4pjZ9I6wdKU22yPFRsn/Mq8mYn6z1kfBpPFh8KjLrW2ml1l7dPCkQDt
BtVDuXWkAGitfSrsVdX6nNkQ6JZAip1WCR9AzuPiYBbEqXRWbMU/LCYH8AS83m8L
QyC0/GEvkI7RS/t8Xa3tykAEQE3OTu+A2Wh5za1LQZcMrj4HlaxVm0HHPwXTD0ab
VApAh0Qc6PXm9BVJrTrGlOAtzXSYNogPA5tk24PIAkf6PcEn6HpV39bCe1xmh9tI
NVOyaODFFwrJt/TKAlibuNxEa1R6HIpyCemPZGnVOcUp2KWXTlap5V1HLbDNjqJK
jDt2EAKrtH9scln2sKsaxXiMfgxLRbjFYmHYg2+MMHwSTRkUm6DP43AjSE6OYfiA
U+HC86edYZ2rm054SREqlfynBRgAfB1+VCLJIiDa0cQY1WBw47p7QZ4ElVO8Hb90
KjPfDUbrYL8AuWcETj09ojEXWs7E1YHtjzV7cUpy/uzOHfJv/vdWWCqDkSs0Zp8k
tcKX9KwA3SFvTS9zskvui3W3vwbssPcuGjvgGFw8AzAtK0YsWXlDm4+u8/GWBaCm
jSHl9D4hWKyA9bwpbMro5Qto5pmYhn5Ow2vMfvKHw1GcJanRfhgtuk58pXIj53HU
6vLWVwlq3t3jZsmCBdQOBa6tLze4QVzIprKG5Iuiai0juAD8g8FgmrElimLqVpJp
GLRt5aqDBUpcK1CtKcgUHoe8u9mbTHgGq7o1zSQu9uFcf6F6iDywgN0kY2dGLPB4
kN2YVGXpjfpzp5rd8ceJ1PuSuPg0lsA2vRW2yv8gQ6ZJLevJ1oX2UqqpKZvM7eR1
4G62ZAGXpl/neM5PFR9eUqvu12KWInibBTV3MoR8s1vSWvVXACefnTgNJXnC/A+2
37dB4LrL49xtOBLUpJOX1EUQpCLQoBfx6eOsHVv9+B1X6oDMIhe7U7fanx/AGtN8
R1Fk4YpDN800HOKJd0un28+xanurUqYdiT064pzU/xLLf1xFFOaQtHh0jpg5l72t
e4ni3T85Lx0sZQw1kl1myLsdgr2/JQ3/tA2n1KnyPi+mNlVt3wUjUV2qncCreoxY
rj9h+aeeFnSrzSLISU/zcU8Ci3eHdbWSzJH1TZ+baQ49OHR0bml3jYlihHp5OSqx
zBCTDFQ3qNWCfqviqsnm4qAwfdgwGK/V4pT4bVvx4KIBNMEwyHxds1rZy6UB8FHj
7e4YeTlMm4nsInF2ywFlnm+uwvLEqB8KI13NHcPHU8M+SUoIRUGj03h+xekHh/KL
+KaZfYWOjqQxyGnhkA+1NbULTPoE9itrjC8IzsJKRf2AbWEJ24fvtiG3egpM5qzI
A+W+2I5uCG6ezCkH2TOgyO9+bRI4Q0xODaZeXxWS+lxyn2gxTL/Xrdxltpqz5AzZ
TBhonThm1taBMlpd+4o8jVXWSxzsypnwrq3360EDm2bavmDY1nNTeLxoM8H6Uh+v
EDT0n5/6vzYQrf1gNSFFDiSe+lWEDkQL0AdmMolaEDmjs0dP1PPqDz071byjPifi
n42D5tgpfCdbuUgNkWFqbEWzleHDKjECyzIz8LObCps3VhF3tRrl+HFw8VrE41w7
YLZRFPmBlaSM3RTihEVd3KuyCCAxYfymX5jEzhJPgHAxCiQGL8Lq4lPFgw02lboq
LV8giJG4NPeRMxQbRtQgMb9hXKMg5RDHJxbSLj0HLnYU3Ry7o+RCrphLDcUx4Zlq
X9BmmWu8nTlzIJdF0AEADEGnnXnAuEMMmBm6HFzfRKwWRd0NyKKDHqmOd3IeWGtj
OgpYDMKhQpm/4GuD0zeenf8JYn4iUm5dxWHC4I+/3WiSzU6Yt7MDDBSdtW/N4YTz
zQ4UH4i7q2sw7hEwJQJECJTSinbN/THOiNQtstMCvNEgVvVB+mvjVqeL+Sf5RWcG
tPvgXiflAWYjuuf0YCcBf549riVXHc0Zyqn02wUFjwc3XFPW+Eo6m4kwpr6XkHNf
9pm+0Mi2TBay3s0Hp3ijd41xAdsKUXDDbvwTz8OFhr2Nw5MsGg0+vdMc1V8hwxpU
jYB0LlK4aAOpJOVdzUcnMIpNmZByCeqAOHZ8HKsC/4Hiht2MlnvPhpeaFUmd9usQ
BaD/WTyVrMfAbUl12gV8PRSmZcplMnmR3osoxdPIbmODm9Vea1OsEcFxNy7PIakY
0dI2WRBGk4vf7EW+CnypCGvV3cWzrypnPgwLS/1b62BzKLVyhFBBkJzEBbwlXZR4
kRYzf4sKt5FH7hAy79ZfrJcmqRemkNd3GiwQjW/8uydFS/UusFsn1Ox6Veq6GiOU
DOhsStkS1BPVZRjr+2WFYbfAy2b9mYqwHo8NGOOAbm66+8PeDPOkizpS6YN5zXof
mcF543pU1JMpY0hjqhMwxNWVlU+cG8+sRAMr2EUq+QgkhV3yolKUkjryzpvixDow
MkAn41nbkQBRcb0f66dyr8kjg3VLIsZYF86l3F8WMEcNjahRujIIu9/DmrosJdYn
126WsnLyuaem7+5EbUeTQCRKzsX52Lm8FCPDUZ3lPopPmcg+k/BCL3BgX5vQqIs9
DIqa9xtm8G6/VccyBP/KVL0+Xj57PuM8FHs57KSbnWVaCNye5eNCWIy+UPNUDo0C
0yatzDwphd9fZ8YBAQu3UxAVYEtNzhuQuZVEcpJRiVtP4/1dFmISwi2OQDT9h9QA
mhdiNR8VoHfYp5DsLJ0uzSnbEXbaFpyBfllCmw+cxf93QSJNn3uTBmJLSYje6VQd
Ppbr6Fqgvc4wn0nMVQqwQ4VqR7RSRW4fP8YLUJ1HAeRGezipg0Xt82YnL39zMnvz
kcLXHT7+P/YYHs3PcfI8R5f/Hy9qWIY7OxiL99swfACX/lo/Iak4cYSG27VkPzwW
d2hQ5b/3VnR4SCbxCbObfHTHNuqmWqb0F7xCGQdktp+TQ0PXKtOf4PJwDYIeQoQF
QVmaw9QfUfrahiST2TBmtZjsbbc6s8eQuMk+HDR4lyEW30KIby/YrYpWXCnqAFGQ
NvMxsV4ici75II3wVmBpvJSzrGHyMIJ2Pml95RtS/ze5N1JYiHt5+GHcQ55Uqx7M
RBjr7GhHAPBHdKrWZDIMJ4apZTkZK2oMerB3Yj95QE1Vr0h6NHqd3Qb415hZAANr
AP0Ys1sCc030rMMwQ7yi/mM7UllXQSNXpKreoIixE3b8Eb4fljgpHfgYrNN7bamR
0X56a9i82mDh/JC4p8HwQ8g082wZTuDKjw4nCK2LT47ApJqQoCAkcUEz131R4qF2
HjR6pyIlriRu/oYFuutq4Tb/TNcrPCa5SSxqvPmiQDlfBqtUaKIpwk06DNEfdYDX
vcVXrGpm5KUv3l6Yf2DL4jqvG4pHHchqLkJXtrCEmyCeOUq/KgnFiNfevkQL5Xj+
Gia24tNXuQr3k+xmvfcI0b67uj0vRWOinc00SrKiSWTFzoQxc8IqbGEtUQb2MrT3
pldD368JTC8F01KeIuT809mzIKjGsjBDytxQKNJSUNxDE31RLhtR05RkzjGEH82C
KBAzsuw/6O9BkfStiS/KjRqUF6OE9DW3+6j1iSbqaYxpCtQxJ1Q9y0JBJP2qRe0x
VHu7nWSyPJwFCPUovcmr3IqZaDqxN1csb6hUfutPzgIJr715zf6r+xUPw21jegWT
OJFxfC7N2cBO9yf93nlnRcsYV4N1rrWpuW0qxAHMfwgIUGBN9+p5CnFc4oYOZPD2
cTiDQCLGGr7KtAY1VV0/DZFXyY/7eglpJGw29+jLH7aPS9nQkco1uJGtsMJMc1le
1xWg9KO1Jitss3UOkHMpEWC7Hs1B5GdGLqve45wMsxTVU8VhnyXV9WLxNzWNUAty
hsWrpVgGmhGY40Ef3cVdRh2EoW0a5wez57PFRYw7VOpDFicQBbxN9WkP5TUCewMJ
IRg4NnHuP1tJzX/dL3cGmnYBac17xFhSQpVVB06TiiVaamWXmQWlmEWi/SDJZlMs
arWP1QZ3y6l7zKH7l5kD/JGahXB3Tl7DikzmYHcL9eSKfnIDqXxI5vs2gbc0Tm84
X+PQY7KRwLC+NN0fhLaV+WasMtueV7hagrdb3OO7JJwJ8bxvJQ8sDPBcXL6qNnOt
qFOJtiUM52x4fAIIEwE8kHmjcG77ro2qbkZ9zoHuLLCmOvZlJ5hPep51LfjvXENr
KtBo0szZXXeGZ4DOpCcyBRYElTxcTSR5H3FKC8L4i+nLBPwJ1EaldP2bntNfh8xu
yH8GBsVpOTSbEZOxUJ6ze2e14JYwodzARi4glxLnBHWv+m4yuA4kSbDtX7VoAQ7M
QK5m/PX72UcinwTqjYDPwjpOemQr8zI1dIk83jSqzwv1ZxNNH/JCrzrAS0Fja73a
7HUHWIhzR2gFBmSlCqSsbXW2EoyRdpfGGblx04PyHcr8scgDM+9Y6jWmYcZxxT8S
fNh1Agz48Vo+WgcMc0r2czW/2mBptIIXSrrIMhN/tfSJfUlDIRUKTCFjeiAXgeKp
PGhlknELVN4QVa3vccUHKCCT/g+OMjFK6MFAKwSNA92HT14ObyveTWShElSu8+GK
ThWfY2hUQg6ieT88+Cx4GbVrKYt9e/rJc3YvST+wHPxH0PhEn71bZj7My+q+xZ+h
36gY3OVduuVNhM6KkzbdwyQWCIvUH6Ehxx0T4S4w/DzyPUFwm5yhSTql1NKsLiwE
B3yrs8rOrnXvgTC9513S6J9QoDn31TxhsnTSoOHgc9yj97pqfJ/J4cX7PKWtHwdU
BJSIzmd7xz5Q/s8tRXAMRzYTYx6u3N7Tk1H1Iv2Kj5EQYm4eJHh4h1EktKFHMuXu
Muj2A4FQf9Dc+PDf7dEFGfRKuvmkqgDIW6usnE0mk9/0e1KBXFynBMzJwSGQ1gl6
WkUiByZnwnbvi0i6rxwUZVWZ8npo65g0uxG9cr3pzdIQM+PLDhXG823RXJ/LsB/L
rN0ksQgHaTzg/zcWdjizOwcVEYgpyMHBoL0JrHix3R0atSHzE2B8eX82viH6XXIK
/WazA2kmLh7CmAz0hp2KU0rIJypNXORN09oCvShDr5+AuJ7nvVnLx1huFQP7KLro
qoJyIAfdOUGwfW8/OByP1kMTMBW1dKBwHTHtI9FiPBZXRWDv7QfyC69FlaNJA6VV
tYKrGYcnYvB/g681DlqhSyraS0WnTScjPeie7u9CRPoP4lgqyIIImFG5wnvglsHh
4QFA0m0DJxnHzFwir74IyiXZzi98mgCu+S8swuxBL9dMg3LMOZ02vKMRemBni/jY
JexLGDFTyWB0Bgb1gj0Ce80hk/naIYZEWy82QowQOLg+jHAfQRA/cRxNmwHX3V3T
72Iu6THvZlDjHVKhdrdsmOIc0JuBGEUW8UX5VcdMVEDAnS5MlOeEKLuHO+Bms+45
cUuNxcWBlJrwVAxwkTouodmpTeAocuXdJDsW4xO0jtCl5FLF4JJAlUxCfOgfWwLG
MPgrYZj+1u8qackFDRc5FEJgYmfijSWWLuGZXKns/5Iz0aW0+rSPN8lc+1hUxGlh
0EoOcmtubHLAj4eFo7ZAIyAboaT9cTUmeqYm8kkXnxYbUAmIOcHH0zd6lRCqKvS/
JkUDldGdc16/3IPJIVopoL2SY/rM4vZyJQUgAoC7jM03B13n3bA2G5WyFazZ0ss6
hUpx7TfD2VtR47OFoXCsL/mal16GKqxY4AksxH1UG5oVhLu5ysJjVnFB50GfArwg
2i0EDBjl9E0l22iM5aZQpqGDqT4EBqGyKDTV6iHRVf223CkiBG0L7yppB7991DIk
/8w1GVwdETA5z3BIUNz3PbmjyhHNpgVRs2dR2vCZ7p6gUocEpmcaFttaa11R6SQi
duXdmRXWMV0MGH2IHvCQv9bHHpEvEJDsRNLfbL07VtaP1SJw1dy6IVNx2QfdoamU
SMp/6Xu6AZcQYrsL+jgYaufGQ30ypEGOGtFwVYBjJYRN+AYX5PtlimyUWYLrTmKF
SmXHSzH82srl/KIxf18vpSEwRQ3Pz6gjIDFkB+yEQLA0OAYNrewJw7/BFElLd8T/
C/B089A8kwQGmUJE5FXF9vRM6/f7YI0JlOSr06mh5/frxFU1Ay2JjBXOO7XY7L9A
dBK2fZYzRRQPW5Cyz101CFKGy34v4bJkAiVskJ4t3CJ1JfVDz//yEDJpTp+TaD13
b2r4qIei6K1BRyVPVkUq1yWMO9R6yVGesXrjxW6zr4jI7WXZN8zivBAfBAGou/mK
4TzboO9dDkpn2UI0WmxFygWf0cc/vprQKsuTMjfzEEkQ0tQqXoPla2zAOs5Cb/UF
I4kdOy/PLBLtaKXBU81IeyJ5KFI+GCINZJEfyFB4v4yQDVuOSjIZqETMApuC5Njk
rINzCwMuhy1v92s3ZYwYAdv/w6e2dgkbI4SJ3swE5Ig8hursEq7HbKDvJA6GxN5y
ICi0LQMuiJkHb4zlnWngNnCItXbHrPBk2sWkLlxphEGymI4CW7zT5FjA9BKj/zux
SukkT+4E7xTimNk458HpBu3qpOOkBMhA+bk/6/WBgvvsAMIVrlF2K826rnWiodWv
G5PbI43aIlxSWmT2BdriuyIqtaQdUTQgdmMgfdv0W5+lv+iZuX+eKVBkqu+kBSnK
9UKcpgZpJXvCTRCv4p87nzmjjzfI4k28CrCbYdSA3FPbEUhywESaSvAAY8eoF+t6
Rr1WLtFSSxmhllXsSw/HdlgkbCaFpGRHL01pXDcymCs5kFRiLSl+Lt1vnSwGKlQB
2YP9LhgCGElxV+HrVpkG88THXpSKzIceNJ3tgCNbV7O88MGh3bfGJsifCau2yYy/
bGYspHwv5cTIHdNAvP0Ym3vQbiiGI5ZrNL4wDTGFYLPV6WKbpDCMxe9Bk31uQkNx
EEo2bHGcL/xymcgwWFKIiJl43bjIcpW3oGsUtYTcOfk9i4znObZgu5Gd8wYyKeIW
Sm48rS3sDSxcpRVAgDwGIs4XRG6RjxVKmRB83STA9v1WAG9Ga0HAWShhrx5p7PKu
r+gn1MQthyP2fl0Xd+VG3tNdCgwTLRmWXciUSHvRwxAwVzt0opH3UoRhMFZc5Ehs
Wmoyu70aozFbasewL4UFKsNurdz5iCroi05LjuSpUNe2lk6zjNtyfbAgvnBmhtMH
ZwhH9iJWDIzSslsyPavtzEOEOSgp/2wQhSydyLl0XmFqy1uCKM2yJr7cxt9IdAcL
GPYnpvbWN3J4iIrGxqpD1kswcwHIww8snGE+JQFsczfsZCEsC1KVdvyh9SBf5wQs
6to1CngkV7+u43Xl1SzZFQ5uAnFDZMAB0R1q+XeV8fMgWBIiPtwc2v7hr2bFVsAn
9KipTaa1NWpJEYxm5mtGvZbgyIknyAOKglAuCT4nr8OdtiXDlWdadsFnBt0VZKVe
CNTtKeCWGXKAfr51RZ8iSYu8TAw+WWT7RlKFBzGRdni8XDTETnjX3j62yMxh6vqI
MrMkbJf2m5YOWKbqEqijRvJXhHQRsPG8Ix9YBmG2tOs8U6sRv1N6IViNRbf12/zk
IVRahmWn55v9kaQgNHD14IWWnOfXNmEQWjdD25OLb1/BDsafxa6VzbXjbVpgHnbu
kgCM9rXpkldMJCmHv4zSsXdj3fLB/Fquq5vNgkCMUS6fLcP+pSseS1MhnwCa0B0L
rnKOFUGq/q5MO66yzqbKmRdB04Refyozr8jAIwMAlOz4/nVJxB6f5moGp0WWo4Cv
0QdlyNmjV8JgsXAio0fy5j4cprUlhbspWWj2ZsxZX7Sqw4iWoAMbK8GF4cgpVgpO
065MU0JD4sGYM55xwhN6fl1E9keSWBG/zQFM5p4uKnTdPj8eKrdfdAUCb270YUpJ
cVO9Ltm4cykxFFVSQVk2vd7QRzqUL9WXw9NImA1P4cGvPjPKkve9q09LZesuGpp1
JjDGAGJzQhAia9nm4Mc029jKem8eFE0A6TJxZWFEdYgbN5SAcTRcyVya+cB91SWJ
UTFyvrl7ntskgXrRHzz7LJHIA7LtNW2tc7H/kn2v458dMFh8Tw49W1wxD6s5rdJG
bsJcHn1tI9gMLBiSqDOrZMGpI0GwsTAqPJrQHVVGfvHf+Igkq7/CVKkScpdstI+0
QlXbMcgkfvIZ7LjisecydqU2551Zq150jy6AVOsSYvgQK9pUxVeaEfDofadanWu5
32kxbm2E+vkIffRaVA7YBpwy20TZ7HNueCulNp0EP7U9JSh6QBhTUcsJrqaWhxHH
y/DHwXg2SMS5RC1UoRIXEQ7eKoh5es0Ez9qRaSrwbF3qS4bRSo9t1a9rQWFb3Gwf
Qleq4/Rws2CBD6nRh4Ta+K//LWaNsTy5d1N0HKjpGNIrkd+aJ1syK4wfC7dFgPnA
lSfXIAIDCE/KmyH0mtQ4ovE6euZQA9yAmB67XAY115eNLw5Cj5Hpk2c34++XbolF
WJ/gV8L5naawe68ioDTU45gQhgrYS+WZp0sjk+2oU/MkYF9QF5Jq44soXkPe4S8J
+z3EHVN4dvOX+BpZZT0P2/DLjMr/jMTMdCwY2zg3uRFAbY2twTKgzPWXpQ8vYdkH
iJdl8E64EnWkdRDQNU8Y0l+jxMTWRR8CHLWhWygLuV4AUOl7owjvA6v2XXYpbtxg
NKC/XIEFHPIEeaRZ99Cx4BtMqZcZK4+21G0uYs16UcXVR2Y+UccAnMcM80/9++W5
sGz1SpH9fhzEogKEIGfXXgFiBxDjeSgnQ1XQHpkvZUevQkswdKVNF57iQG7cjcgB
7sIbhzJpFa46Unvsv6dINA4AVnc1gSd4Ks0yQel5LQxhSZ5T10feTGtdcvEbTAWz
629LsBYurkpuVil6OvTi1Kma1PwygkfAx6I9DHVlgdjxMlBs648wxyPz+SpxTKnZ
aBf8A1LtbBQ8pfP3e6A2RN4YHDWRKymZv1sk30AhYzTd/2OrCIBFjEPzdEZXhe0N
oU+ZmNklECNJP3pnOa3B8gh9ym/fbcNjKrqtCn7L8kstCO0lYOcoS0gHUbvFADzJ
gbsZNx5H72y4EO1u5+u/VG2kzpCo+/7VOh50TkNTiEA3dAqkDHqnDnuMqtJHOk+N
HiRAylq67Be7/7K1zR0NOBaQmhZcMyjBBR8gwaiUM3R6ubMGTpi+ByY1P48ru0d6
fHC8Ud5UZY0toeIyrDXSoKAp2hilQYR36Md41BzReo/ZRnNyElWGvSX7Io9P8eRb
MWHvHMolVWHenFCCyHrXar42NpITV3M5ffGjNEXCdVtBYzl0K9CAqdci+NDOjAiQ
u0bLxFb0c7hq/joLb4Cry//DfmX56dl/jjfliwNwI1jrFmY+2Vod/QTWN3dUkt/r
yMv5DpWfQ31leHgS5P8HADONW5VIrFVmn3CcYsElJnKuHCUBe8fjMc2VJswyfW06
gQXIbvROlRIFErmaAaKQ/gWMm4XNzxscKugK2fcNOC7EBn3ciqyerbyuPGPwgOx2
PFn8iTI6PZO0BVo9qiaINpRUxbZ1bvxCmzcx3wVWoxRJv1dM9RHlmEsFhDfB63rK
vgHGaI0TyohrqYSIoHDcm8XC5hahksFl1eoNYDBbNxvrXjHFYvv+q7lgSzkpRX5V
KTylbe3WRVU+b0ngkKc8RwPGA0NMjRAOYGqtaLzjgfW90/QMGl4dn4dou+xPqO9M
8qg3boh11uVpKf8/duKBjI3Yad7a4lb1lR0FIHd+mElvhC5yuth6m6TVaysKoVnb
n8htTwLTK+Ip/PVTo+vzS1Zad8x1KeNIBwBajv2pqKDbd/JVw4qlfTDA9WYVpQ1E
7tEQyWQ411/hEIyHEYMPDyx/ncWoQhxQil5iWkO1uL1XZL+eWPJaNxd5VMDVeF/p
1LxUXtEUIewM50dLLbLxDRJX2Cw4s0n7ye3DQz1PI60zxNDptptMdoa1b++dH241
ZBx/BJM9c/OUL2ogpl5w61QlEmRZI/nIai/zLBCEyvfRccOd6wGCqIO1Tyu4lG3d
P8f9Yf641rjv6QxToIIo4aK9A4MJOWy1C8vJNSASZ+NHsRPpwz3uRySSQIEmNHnO
caMaOZiLVylMIilbB5BdcmqPlnIgIKkAYZ2WQn06xPp6DBhCLI9HOvVNK9VxhPb7
A/QCRAK2y2xQk7TWDzs1pRsDidKVCBUUf8ddlQHr11U7giKGChr/ysv3HbYf/4Iu
3afHTafLslzBJWJLoD+Lasv+zWI9QFkc6vsvkuJGGLowX8GQfXQSkR7drh8wZyMi
gMzEi9IKAK4TT8JHQwuFMZiMjMqMrEIhEa6v2QvrASattHaNIsQhCq6b8obj2CKS
ruOlVTXo+oIwGu05vHYY0CiBYiLWL3sMUYqVF59nbHdLyqSGp7+UB7fgQuqpWPWK
kMAraT6bz1V4orlWuoFWRE9bMP/JB0sWnV2ZxZwDQRqCTCYQgVR+K+AGyIVh9V9L
SLdNxz3CJA5b0tAuhwHIFCGK76FDATwhRkH1ya+AWEVhGUMjlfOebxSRakTSh2cz
U6zWpbCLUMRMCl0LbX9kRaRMHaPIubHVYKQ1qa8CdmAjg49xTKosEprY8YPGlX3M
M4J/KOgwDPn1kirxr7v1lS5gKOKUvPtbdVwyNpH8QbBvhLsivtCkBrK6RqFUXC7e
z2CqKxKBY2G7Yi7z333iws79sMhmgmvp7rKPJFyEMK4wnDVU4+V8j74DtBygRC/T
I01b97xLvYCi3dtj8hluoRw9paUPwiBj2tcPSjXfBHAbHwAMgyYLKs/GQQTYYkIu
6zudgoz7w4KkdkMN9cqz4IeCNg1B8tutRRfUkc96MThM7/KUUrMiy4a54eGRUc07
mGCL/kPDva18mIA5AcPUEvh6pbRcz7VbSdkCPcDaVaJ85g1GmFQoB7iPj46xRnDa
mSSwsgb59sJdzwz0Csjel+Az5P6OfNEsdRHq9I17e37fWzORnEakzIPd+adefXFj
N1nuMrp04+6pDZ3z7RfJSvhnu9vOgHheTJvvStuu/IYH8rOQ+4KVY1j2arvNN8Di
6hgC6Gtb4NCoKCQo53WbVTjoycwg7UJQoHgGo1DiLHci4cYUb5MTMuegkRp4JE97
kHbb8g1A5qIWiCxw4KOsA3oZA2uKhn4ZAC232Wc39Nj7CQYXUqucSjJhUjeS42fT
BsGSmTd7/mVGiQZBSAxasODWXYCfPtJ38vaOoot9pXqCDEhmuJE0VcZ2nEn0rW4D
9OP82FiHpIdwhVA1ZW8H7FMEoYIrHRoH3qURFtOWvtP0qPYKmYvajwwh5v8kFO45
3LnleYYMhaTBJxmy0yoYqg==
//pragma protect end_data_block
//pragma protect digest_block
M/BAOkK4S/jjAzE4lQAn7IRMS88=
//pragma protect end_digest_block
//pragma protect end_protected
