`include "Usertype.sv"

module Checker(input clk, INF.CHECKER inf);

`protected
a(/f+1cXOcJ]7;V3,W]C?8HdVO(6+X1c-<T:L>D9YCg_3K@W+#\[4)4\<2bQFM20
1X,VbcF=SM?Vfd_.(?S]_7Eeb02:5P/Nce\e<5;5PX##]J)I#5JHYc.+>T5UMOGC
Y8^1TK0fXfb7Q=O9IXd>7]YRA^@BKW:S52NSA.fDOPeXPgI^.M6M\=Q>)@)K=F<O
>X?DgTaY,bV1G_(OZO-;]dR)^#ME=?->gK0:Z)=K[<6&<G]JbZ<TE=64M^@#E)SI
g;SG)^HKRF5PaYONK7-6]^?=,8[>M.e#P(AVE;TBWO.<;TPG+4-JUVCY46WWZ4YR
KdcY00MZA,?MHE8?c<0I#K//D[PM[E6.[:JXc-[H#AOVLB^Rd.+F&I\FL3K+3aUL
,a)6RT6:N\CWAd5/LD:AD,(+R7);Q=VDgIX[J>_TARI7KUSS,F,KC[AJZHR=[IK.
+V3fEXN#PM/8@T@>&BQbYR\C:_:VC2^4_=7),NbR0Z:7>^MV,C=-DO&.#4g\dF]I
MD:2[^../bK)HH^<T&F=&N.eVT#Wfg0MD0AU3.P2B)cR]TE8U9;aG-;U9e(3Fb+=
e8YUYR?Hcc8Ag7/I?JK6<FN<Mc[2;;Z@\9-eg,-(;NfHH56V7g&b2UBI2#ad@RK,
7XC;/[\53EH>K\<MT#J&K[^:5BJ\b[?2FJ:J0f-AK<ML\K&d1<,X7]IDN-S^1b.4
UHRS=O;e\?=,7\.Tc)MA&_c4eZ-6AH5;T=g_&LXP\cH.7cf:70;B9@I);WCgR+A[
=RC/(7#ISg^ZZ8.H48FQQ1cCB33]Ua+L9T;6IOA2)gP8Ya:KI<O==QD]c-?81g.Z
Q5[SIP-O7e+E;>-[DX52T4HT?/Y-G#YU+T<P=W64-fF_MaebX<e;K2g-e/G+1;SD
.LR8U]YbbR4[0_WKc-V)-@UO1.?gcKb334aPTca;[&M,DV9W-;O0=PKKLDM=J\D9
C-/VU^Ef&P0QWD_SN(\g/M>T1)ObC<TT_WV:f.708EDbZ._;>20G+V42aM4ebA^J
)(OcdeO^>_?DHB?Y:_=U^#_&03VHR3MK61/#?9V_D8Y@=(gV\,/YG7GD&8D5T9_-
V08@c,WWE?NFDTDaR:(XZEW2g6aM>U6g6MNDJWIY9SYL93KB>d8W<S<O?0KC:TSJ
015+@#<#\5aP5fcB<&=7XfKKS\@c-Kg@YPXWY+;=FR=e\&?6MgSG_MID&:+FUa2g
;EXaIc,4^XLD6IR(W19c:BgU,(TM>cUb()d)9RM?0)_)J]I[M;[0B27_NBLS6>8I
KKTC/gH1JJ<33XYY6HGd<.Q8</cEeMWBf&VQ).A1O6gR5>.7C]G.S:X0<H7JRd^F
K4X<3DFU:R+fO3,JE;d741X(WSJ5ZbJ?PdSWd+S=\AH;Z&2GD87HeP77JVCN,GW(
XX34gXR0+1A6[]Y]X:UGbSUFD=HgG(\?/65c)-4+G^d-Z\C3?a<D=Lb95LY[N#Hg
LX3>4Od6HA#d<&ee2M)cM;[5/c,WfgbAb:>\E=(5K(A&<EO6@SB24N/V5_2S^VGC
:JM?C(3CIWMKYQDMSb>XOMR9_AL^PZeMIKg4PGaH\eH_+I6A?QZb[+X5N_;[afa0
AI,HHZ5Oc3O?>]RVR+_D@;97Q<2MJ;aP14(@NeD[SB\Te>S@Z65;1Uef#H9GG,aW
AbW9EPfEg@e2;_;BW1JC.IIcJ[:H+]Ge939ePI80H@U_FGZ(FO3?>IK;W&UGdOLM
9bTc^2ETSR8VQY_KGUW7TQf##QP57],KgRW8N[X?Xd?JH(3V_Y[^7efAXKbg10AC
DYGD(_eH0>P^-[WG;gDWEH:HFCAZ]F]UNYP@0SLLWEBG<daG-2P,Fad=aF4cOZ4W
bD\\5d.=+E.&XBY;\&?>G.3PJ,-OS;GKgb]8Ye\LU@=2C:d&APZe^@PFOb#KGR2V
c)I^N^b34L3:g_,-&Sg65c55d=A+UIV?aTPg7KSF8CR5dN+S;X+-RTZ80Q^6#=Q\
T\,+)4\3L7dUe,M40&7GPXf.+D2_Q2\6&\N&[]6Hb[3:B8)GDJ7O5>-7D(e<3]UY
_SVa#^.=YD,R4)3POQKb]_][BX@VDV=\TO#V@K#:9WW\JTCcfY4UbQN1+R&KK7SO
c/&Jg8>KVa,g4.M+66#6_S@M6RW-c@G.#6\RX<\JFCM85(BM>Z(e1-@IgL3DHbCa
YVK:PEfc4Tb_K2aaME-Z4LC@DJ4NV7f_JBCGF]6f;LKL:\,_X=0U?&ce9QIC;MLf
fG<FOaEOM=7BGf&f>3gf?I9;TO[cDNSS[Ea_e33^e-+,BN9GB[F,7D_X:Yc0/Rf=
).CRYVFVR0Q]BCb=KRD9Wegc4]HU(a:XSM[FXLDIXYVZ83DY&;9@[)&H.g2aYH>E
X)E],60TYV,X\?MB+M[.K&CaOOa1D7>C[_g.-fJ0e3E.0g\DS,4:D8F](MNH/&)[
IJKg@K<BR.X6=1+8aHK(c4e=BFQ@.M..c;@S0?Aa1L9KZ_P>D=c3K6,9ICURU#\9
OfHb#8P/\46Q&7;_GP>V4MQ,OM<RYB[,7E+,B?A-V/?5)YC]R26A=@6QNFg]#TL@
Af_=V6[I@e6[+&6UU8/ccg>59&=71/3)D@3bf^V_dYA;>,ZI>AJ3[a;(_S=[NgKV
0ZR/6J_VLg+__/Rf,[.SQ<TaF8WT@?G@a)/e1]1M?5f,.9e&313U5QO-KMZK>;=7
6_5N_UO]=Ag1.ddIGWGL8aBKPTaV-1XfU&50#&VWIP/fM6FQS/eLTZFL#/:Yb/5U
U]A7_b.)c,]5S/CaWY^b#a6QH=R;PG_G6CFNG;fI-\F]P1AM,I,Q&bKZ2/9&4f-R
.9U=Oge,-,8XT\<0HIgFRWI_@J:AP.\K_UU=#&<OR3BBAXeL\7O3c[SbHc@?B?T8
N^YgB^]:BM67#>:TB/74OD/c,-91P1[[83cJ3;U,5^+Y6S,IDUJHVN+7YGL_#aGD
N-H-XBH54T0=<5+U6]BSES\Q6=W7<I-0cJW/([a\a(8<SgCH<:-0:\fM;JGefHD;
V3J.NDJT=X7)a[CK^@>;D#_).8S/RRgBEHF.DU802eZ;G>,L@P:;(;3/HZK[L1fd
9IH/&]gNJ/@U7P;69eEYdB1d/)PUVg#A:+Ab92IA@GW6?]OG@@LX[5#V=<N2_ag8
,KF0?5W1(gg+K()(CD0FH2._Ec0-D++BR7,DUe.;R7eJ7>,W^XU>U4\M<3>9JA=0
S#,>K+=b86F0<JZ0XXDV8:7S.JT>dRDC[<X=17]83@F9Y36##TAG456.&\Y0.K]4
.f=KX6\VFRE_9V__B/BWe&Da\fM[-G71M,<^U3@7,5V^VeX_UTK>d-&OKK8UE@L<
&5Q_[cX[9^bE7,W<C,7dL@:B37VM3321)>>e4F[f_@Wg^D^W2_@#9V3P(T:N\273
/:JeO5);Eb9Q-ASNc]7VRMU\MQ.]aHDH9d7\RW,fZLf^?3[M-=&/<-(W=E^1N7Z6
&NNA#bKgJBO3#.2>W[1KG3PH&IZT/8NLc^f4B>1;bfA7G68bc1EO4T\3/WH(g<C;
Q1M)2]3CO<e\6GCSTgN96]a/#2,V-,FY,&&:162bJ&3EMUZ6e\+,_QBQEa>#B1[)
N77J+7:&=F.Ld+:,fLAM[[PL\)IXQAGeME6g0MU<R0K28e20?O5.,N/KW6Zb.@&5
4^-.+@:PD(4=(Z/7AfKbLI=-YN_Cf0BMfRQ_0Qe:dfg(7K3Z[?M1G7MfWB^cZ6D)
MF+fFK934MD>1HS.5EeGH4RTB4(9fceILAW.+-DDDG5RdN,#JFI6WA6?HPd.:9>d
LRSKJJ#;?<AfCCO@c>OA&T3D(.S/V6A9(;RHAaEPI4],D^8[W+,>QVcL3W1[MHH5
00OW@2VF]f;TI[K6835?0-_eO#J9GHWD70>[&+,gI2Q80#V7FTJ/0R[2bV,S&6D)
.6>a9bO=G8=Y&58BZD#0_X1,BFX-X-S>3:9URR6UP5@/;fMW41&)+ZUA</EV0KL,
F2\(VTL90<Z7TSIESZ7DGN+6V/<dGZLO]8+Sd_=^O@#[9(<-MgA6bSSbY&3d7X0=
Ae;N&JWCUg3J4eX.#X@QFVEX@):g[b@PB_Y/Gae>eZS.THOL1gH5bbW<-d066]LE
6KDL?ZfCUCH#b5G,08=.Q60@VY:X[YdAd#Gg>)gZII>?\CS>eJRKTV:5GT0XO.RI
HFXNRUE&egL[QU/0H0fg8gLDU?/D;AWV77Kd38OL>VT,NDTgPF85aeW:;:]ceP^F
=([]JE/TAUVgf#7e9:0Y46E3K_e+8_0>(?LFJS2d,SX7N9DZ6J@2f:;MU1N8XH+e
[=ST89Y0[\:g?7,WR\b&/BA\2EW7E@P8]T7-U[<@S<Q#DUT\#d9?9H]8A>KB741D
?\C_#&10FQ#A<-OY1&Y.V(A?9A]SE@F<G@.39P5fL4A-OMC3Q2?<-KABMGe791c+
UOb)a3(]^JO?@0XPYTF>V]JG>5YX=eB0JPDC(OGP\Ca-2-2)<YP==aG/L3V:LKgR
CB\]_>CLA<f@.SYVIG@3c_8(CfW:H]6[8JJ3?eXXI+5=.#NaP59YH][WC)RRcANF
Of5gZ8,V;g\809EKOX>U]#2II2[>Y1AO>8D1&+F,2)KN8?63B0Df.:0Q_I(S#AQK
^BN1C1GZI-I:b^(A\X6M&O\SdWKf:B^_d0L9d]2&DZ,N(<2[N;OJ13VQ,O^:1gZQ
YN<E9A(:7_)E?CWI1DQ]0YTJSO&OFP5&QAV;S&QC;]dINeV^L,b\F+cVXTG8^3,3
A)aO:@UcX4YB>HKXK^SLXH8PPKUSY^fJ2I^3fYfS2;4]0]7]Y36(-2ZSVR7>aS>6
OJ._QK7(M9;C55EY6Nb9YJN_7N0-JMS]KdDM56@;Yab+2Q]]E@A^RGW/CMP0gKL#
MZeAeCe9C\)>+G^;POaF./<d@#/fYG]faH3HT[W7/_MU56WCM=&:_H=X58XY7CLC
M]\bL/,a:)R2BP(X<)#,=eS-MG1g,/Y\4W^PX=&JO\a>QA-CORWX2U):HfNbSGU<
UgaBV;.8\91(1aO,?OLM>.JB]1fXN9&>:&FMHGD92M2W1(P29^EgC4g@eIDJ5EaD
YAYF&:.^?;<^D_MBPWd4e@Q0E6;JBfWQH&T+A@a1>2NJALf\72dN3(a&?^D>WeOR
,-\0B\T4OH0;;YT9XW0M&=cdU2N-)GISJKg^-LNSS=;fQRT<BR2a]OJ1OJO]b8.^
GKNc>f?XXa:PH=9Z;cJQZ8;9e+4MYe>B0,?9)^a7:X]+,;a,H]g+7H]QY<[Bc-+\
FD#)T@S:-4g08(dPV[LI<IVMR2&<HV-26(9]G:O17QL-R\-bP=7,3EH:1.[-91fE
#;e#d,KAH,:^VRL,[Q_5RARCM(3L]f0V_&g5<H^YG6A]/?H)7_DGb:+-04IJJ@?g
SP^JTJ10HF)=@2[P=Q=IUfEcO>Eg[d<EAFR#>SA_1O,5\#<JW1\We1K&1a_)FRJ,
d6Z9ON@GV,G>J7Gc<B7J@E067VTZD->HJE9a=(,1FAZN:0K74ZWAA(]M2CVcWc(H
Jde0V<&2)OQ^^72C?g_@0C44<TOc<[)L6WBSGg0_G-_-=KABG]c#0g7K(K9DDbFM
8SE\CO)8b;dZRY#dJbbM,g-0>P2XX/NTN.Q/NUcB\VXQHA]-[B2I@:SeM@^W@eWH
#EC3C-NSfHT&65EeeB=-AY<bDL\\]:LE>NZIJU7f.\FSIBHQT6M#EZ]K#_R-,4#5
/39F>NdXB#?M][(SP^aC#U3^d^4:B>dF6Q8P\.61?S?ZQ]d8M,;DbC,?1O\?(ZOF
5ad=O4g03(+BEK&,\S<N?Z(1=H8aSBV4K2=[,+=+,OW@>?B-F:6B_<f^Y,)MdI>c
>R3:+O5W+HJ-?1WQfABWJ1aXS;_db>W4W2R,/E3CU5+7-FLS,(:RS6^M+(^0g5(F
A_CXM4C40.\P5WPf)<:[12N<DS3PTgTQ0K/U3@c6FHL=_A:MN(aAaW)G13RH[[.P
M#\YWW@TMc17+N,5^?V^&&3]?N3&8QV4&E15H2,^?JA=>O@HCU4P<17K=UM;(4&-
f2-^3^SWV1L@U^G.5><3U;48YD7bQ_0<0aRFNaBZWM+QH0+d.bK3/LDdZf?R8IT+
N7,XBP,de,X/U[)?(@J+BF2KNCb3E03,XJf2[B7?gR7FP38Oaa.#&4>WE7V5QDe:
YG:C_7G9e]/K[G;HICBYNC,>M/Eg6gV1&@-4/R:OPZe3W_1QDbQ=dK>#Ub<@U0<\
VB#1-1HIC^)IHA?g3@:-]6/S56;P3IOeYU/gRG\dgV-)beRfO(<(K5P[SU6:N3IR
,[CQY2K>K6Q4:RK7?E_\6eYVMgCYQG5/9e3cA?/]b-gKN7O)-f_6RPMM&7E@a,6J
>FOP(5I9-B>TWf1JbX<:f&PMU,KGdS##IW;B(3]2=FBXBRKF)^_CT47&-M\4+M(K
/SgOdaPbXT_,]UNM)fHP4U#PMX<W?_c-1=ed@,OWc1a1cZ:HB2XVa9C?P)SSI@c>
H2&82(VOC>MFdT#@M8UT8/O&#DcVG7(41Y1\43LGVZLd0WM(7E[5L=M<(FfL(8BV
6X3-[1S(c&g8L8g>4.aU9=YI9:ca#^.^b<fR1F5\GU(C]J\5WC7[4b<0Ya?X4TZ9
>HBQYGe=7d;8C>>0.a-ZR^:J8C<_?LM92606ca/+/Ee-UZa=8L-eS?fK7RWX.7?1
<cf\)\KTJQ572RX1#Q3.J#/+C;a4.)Q,V>+7H-fUP+2]24b#Y<LVI89c04G2^4Q]
&HD2;AD-U8=?I9O^f]9MO[[7g;PBO:AE>bb=5;84/K+DU]=^=290GOgASVeCJDCB
LQ_ZC.D9ISfcZ5]S#ePdP\RTZQ16O[(R^f;&QG0O=TK??M(\YcSCLcXC?)_M422(
OG:DS/&LF@dLeDZSM3U:Qab=S?A09M(35_F5(K6:D.LT9E1UM6dDKY06.g5V@[#@
aE=K49M]7;D>XWJ#D4C-^>aeHe&.787@[2L[cDU_NNfg9):7R5fCaX8G_#YL+WOS
PdN8,]1\6Z.:eQBQQD&)DOI8=4+HfG>6&PVQ1:#7SFH-C,4fbf1=&W>(]UZA3KG<
HJXY0GK9M5X24KD@QadC@23\ZD<4TS7&<M(7LMF_B3@NX>AbBfLTJMNEe5AI7BU_
<_.>b[&5#U+LgYb__17=7=DVL0;[+0^KK>1XPPST[54+U1]LbfDRJWB>:/APTI#&
;;\U3\BEb48KgX=X7O4@^;Kc9[QScCVW#+@BGd#FQ8.X[-08OJc8CO]-Ub0Oe;U0
]+@LE^-Z27e&OVN[:6JC@9QMHH@?.Hc9_;ZF#c+6.6XSE:.3Y5f[V19N,\<V,KE-
WOGNU>:+Ufc08P@Z6XK.A,:UMN>7AcRP66\[#1Z;a?Q@E<KdEBL&\g+TVM>,FVLS
]X@JKY\@S>N-2RW#P=gRWM1=3Z+31;FQ^c[4A0V=I2/Jg@R9=&MHKLc1JEPG=V(U
_IbY(:51,D)W7DTFRF6JdNR-aN9MKMe@VH&\dc/cY>^FV9_E^7;JS[-S>:H+<S9Y
;7UX.4cb4B)1bI6=J]47T;b9e8D[T,bR=?Yc\.ea\@FLc&?FW;+f/YZ@2g?gd]W)
S&KPSOF?c36XeA&aK2@)TK#^b?RS_1_JT<(R:c5g?NgV;-=Ve>722=0D_N@+eXF5
:L)&eJ+DKP-<BKa5c2];VE[?^I:LW467C=?4#d._E??9EEee_QV)8LN0Oe0+<]DB
UE-IdN1.&;#5@S)4X^2.])G[D2,,UG04gb7\A074PBPUJ8WH\(>;Q?=J.QLHDCdf
)P5>c\NIG?MAM9.?9IaCOVNd&JXR>DKNU#V:A2gA=Y2H32S@E#9#eYEUK<,+gc,E
c.@8PaM/&<GQFJ]8TSDE1@E79]9)Z(DN)IBRQb(L1YOgUWM:A4WQQe2;U-<<a=\G
.^G[[AAf]HA++B2+ce><)/fXCAS^)R)g/QLfD:@P>IEO)aA0CJJdK+bK?9<Z4^;O
+b5c/>C4:LEba;:;.6N-^Tf=:[OG:0#\aHU7_>afVB628?G_?EGVT(0XV]TagI9+
PQ[70gcF87OR(BVDY4;dUI2QWd?C[U5P95,?E<5/UQfJQZ]4I9W#:S:fbP?HZZ^)
>=(,[@<+2_:]cBQN[.+UOCR]X6bZJW.[DGbE#CVa7UA9^3KYHXK2P^.-^:#bC3Nc
e6OG,cQT(fVAAIa[1FJ?TRd;U.6[2X6L&)5S7Z5PI2)ROI<?c2\RNUPOAQYSKUI.
>-1:=aFf<Q,YP^_(1;[_+2R,1^6HO[D=O_H4=J-9:Ia5eSYK><I5\#;0WLH[.Qa]
XGM;/_^cBfbE@14CLV0D<&gUQ=PBX#eb4-44dMKRU^RWE@-ANcYD(0RXA/_DRG):
\+SQI(eL];a@MKRaGN9[,RHHNZ+BbTM/#UHH:ANHR@@e2NZ7e_04+F=/SOUeS8XC
YRdaHLcaW:\c87;S:8^Z&]0FXM/0f4P(LFR&8XR+=e=J,H3gK?fR#D/5FT>55O?Y
/3.DZ8TFMJ83<Y5^SGDR\4>P[#fU9OWcYWc+bZa&OU1VcRPY&g\LP1S-E5<28JK&
I0#>(^K2BVA<JH<b&AYg2Nb;NQ(1T]K0SYKC2AR2_U)HLAH\ZIc_VOF?CBTTP-45
<-U/FZ8OIWHd<P:G5996bVZ\>+2J)FZ#IG9^@FVRM[cJSQ5+G_&Ee#&8K?NF0b3[
UHLC)&--\>dB)QcM^[6O=-(ETeRJa(WH)(ZbSA#,ES#E/HW8AF3Pa1=N6\F0+/>B
EXRDB:RII\IVPae5-4;AE4Hf9/VGKIU=f9T=P)CCc8XcB(:ZK,47]I=0V0QFP(F=
WFL(=OOOggLbb<-\bF\;ceGSYAdZRRG7&aWU.E\E>2U-SW0S:.RBPS@3f_B^DAY3
O3dK3>H;FUaCfD?C<R&3[\F+B:-eF-WH^S,ITXf#\:AQIJ?Bf3(7:bIW(3>.G/Ce
N4?Xe;[Pe.9(LF@d6/85KGGM[Nb.d7N)C\WXM8+;;+:)>(7CJWaQD)09Y:NL;80,
:>:UQHS6WcR@;R3J]2S9=VS+?;7F^#1<76=1:\:&3?X\71NB:9gY2/NIG(FL0FHL
e.2;4G02Z]\aUJG)UJ7-<c5)f<f)eO)WNa=Z-Ef&-Ye)a1@C)L3I6M8MTJ5,K?\-
.3Ib9d&>aQZ(O7?PGC_cI^OY\Q8]D[><>@cY^bT58M.9T/=(),2<g,>O+P8>^[D?
1ggggJTE<_d4+V\JYA]CI>4EKLf<aJ:Y=84Y]>E7.9fAedW@_7N#U);?]ND6471E
A(g\N-:0aJM&P]=E3)INU;a(@GJ9L>ET<>YDL?MM7B7G78c_f#5)93^?.V?:9)bZ
D7\W+9cR1gdU:Xf+EA<Ace-:JL-DJ6M^RBA-#XZ#-K=&c)0JD517RSC.1C_WdIa?
bL?f/RYL>Y02EMSgQD)>]?7>WN<LDH_/;)M09N5eQ^SO=?gA_?GeFT,XeJEIR,J^
W<gZf&4,X(+5PW4>bB@89d&c#Ca94-KE0KV8=FEWCGI2f#0-/Q-SV1,^P9PD,0S(
g-TgceNM25,J>?RHZU=bH2U.7O3H\Kf+Z>8(5AQeDSJ7UKPCe>1BXV.W&O??7d\[
2P,6P<.PNXA5>(80d\[_2A2bGDF<F7^57MI90YU?FOD5@6,LgNI=\cQEUU8d\->U
;W1M\N,R_/Z[DedI3RA=K>09]JNV,8-O_Qa7V-SI^J#D#fA5B:IfTGTLG]FJYdWP
=D52RB^ZBLOVf52^8_L(gW@Kc1:VeFG22]<4))2A])]T#PHK_9e,=DZCC#OF\/aG
20SC,OKQXIVP-3@^]\\XV2Z48BHbcY7=#KAKeSAVMK+GE;B:bH[/==^&(>FOCMT/
)N_b59Fc__Y0A:gd^,Y9,8S9A5=UE2;G_GN=(ERR@T_-#/X?@7f\Mab3M/Qa[38\
beK:NZT5CG4A)5+W[IT@&:T]b>>g(^[K&<,?S-W9U7TJ@1YOgP:=V<YC>Uc+L-<9
a5Id\TR#GZV_2E7e?@0?I0)(&,^+df\>3[FR\#d^T-A]Jd+,KVXFb^=gF6RBU,4@
-5J.>P@IJTUE/E>S^g7U=^^265G,G6?V0Ng9DA29Eg4aGPLIP:88L\LD;?(b[TZ+
#bb\XMQ?O^8+T)\cIKK7&7fL<gTe@XG<_\/KP#ff2XQN8^6MZDc/8Z>a42L_E=XN
@>8US-gQXffL]QDTU4^-YYBI0EEdIg57\A,K7NMRL-9.Z4NRQ[e3cXKdGa;;0aHR
-(&/N7T?c-FfbdEQ-67Zd/3&g?Id>1Cg[HU>D7(]SWYMPH@g>=1AMSWN=ce<E)_L
cRedP/6OJB,WT.&P<,4DVIL>J+T;IJPf6,Sd[T?YN0GSSGCYS5[+[3??+d[MZ36L
cEH(B^[6JB_HT=g+YZ-8<48(8MC^aW2>0((>Xb^NQ,[ed^N)B1(5d9&gcOTZXR[_
^X.cW5(SW+&IfVSGAYeDd@W83CfL4Z,8J>W9VZNLG)Y7T/cg<dB7(@:9;RYE\(^J
KO-[=6;7^f-TBB;9g@.b)2J8/Y9NC)[).dBFfB?/BNb;(M.J9W@G:?E?P((CF94_
/1YOeD@I4H[6\_)P<FLK,+85ZE0[9&g:a6VZW1W(36+B(g.5>:Z_L)]AXbfGegMB
(WO5aMU]E1Wc9:JETgF8FH9N7V[(9\N-(,AB;?NbZMN&>V82QF_\EYDKbC:1c@&F
OZ)OTd^Q#8YNLeCXD^T+47KHC)8IL5KCPZQA:S2L6Q\^VLd5?A+)?c[ZH;W81?D3
+D2ScJ;7#B2fc7aXP@PE,\@\^1_cG=ef[X>AMI&+X/&2U_dDYXZH3^?(A_CdWZHe
DB5;L_X=U^Z\A9#b=9KCE[DUg((/<MAEH;[EY-g#9OM)([0d@CE2Gb\>aN_06N]5
bY8g2&Y.7F-A[N.>cLIXgb#MZcX:b4T)@Y.c#CQ=>bE4aDc8.PZe^?\gBE+]GNPR
-<]+H7H.+?3&:##+):\FcCM2\fUdUQ8YBW_eD5UQQ:B0W@fAVY\e;a/(6g/G34B9
A[Fd>/,DEJdFH9VQ&6+LX#b>1-[NeCfF2V?H3ORR#K:V+JN+c;_U<)?eU4X=&K\S
\.UQ?==IS_g:S.TJTXY>YQ5a[QX-OLKfb/I=ZLGIX&VQ0NMVE?2Ec=SfAcCH@Q]K
-B-cA2abafb#6g6>=0^HD&@N-^\43)Z=c7#AWgd2)=#M.=RYYRb[TBQf-f#(@cD=
:X>#F=g8?[9@2&H4,44S_9A7JF>]?+EO7H:=,Se>LHJ:36MU&JG8+(LPWPB7K/U4
?AZ\IA-G_LfGRAYa>R^^:a,2C^PJ+.M=>UA7=1\OKNP#K-,1]-])8<aI,P0e=TI2
_7D3g?DN0YTCa\+3Z>/Q8[Z:=V\<,fVS&eJa=;:EYC\C?KW1NT3dC3OUe:ZLM&BC
+_H35.#+R\K95Jb-3MUa=G-RI;YM;(WP+cW6[^L1+&Q_AF.J]EYe2JY(,7YE:bcX
-_]AWJXOQKB&_J=DDOYQcTO&e,YJ]J]KQG=[B+-NVCC?.T2U]19/8+@O3;)Tc^+;
1HIGa-eDVO,#NH<&=L^SF/(^5U.ZC8=9aOXeCHYKBE6d:.4C]gH108E/N+=:Ze-E
6Xa0-X>OHYM1[T__@5^Q.0WH?_,(KWQ[L+Y,W-9ER#K_0NB86<U1IONdcGPfD2^a
WK2#2XHG0M>PRPC4d\_bg@8e;LKcW,QK>)GU:P<7R49Z6d-H<LMP5JN<eZ5F(+F[
dK55_7Q3,=:aOJ2BSM-Ze,^WD9SQ(UJA-G-@-1g?,_@N7##ITf6KG1E[]7+A&X)C
fR<P#--&B-a-O1B?Za7Of>DJcM_40^bd<?NN2TFJ6e>4UX?4[F[gI6P>NSXU3\96
:dS;eW8gWHG+&XO&3JN(NPeE:9F^Ea:EKc-gG)=94XJVF^1F&f@D[1_dQe1+T]^@
X0/=L>?bAQ=VW13_e[?_3cH@V&Q@[O37_AMS/M+G-\,a@&3W/ePTR2T\e/:P+1:#
KWZXSNMVfd8_6332ZO,TCX_&D3)SDaV&TKTK13Y.LGb-SKO_BP9I:\L;KYA1O;3O
/Xe-<PTY4Dc_?&58QAJ[V<JO,DF?4]E0W<_?16d33@]=)X>R60_d9ADIbP]f7@eW
WCOJ@c/d40>IDJ]=df.g0U69,a@)A)4dS(+b51>b#.T?X\B9_M-WG]9+-NG_]^+4
??b6;Bg3K:W8TI4UOB+-?2Lc)3+18fZ+F,We>CMG-MLMI1J@fDNcT-3^[INf;cL.
>.N_QXO;+75LFAaf-58433\.FY,IYgZLb+YR5BY9^(6,R)@S#:/5<],K7W,1eIH2
XK49/H<V@96)]N-EOC,V2g7S-CQ5eF4bQ)X(VOB5HI8Dd7X+D,5[TUWWJ<ASeD9R
5EfIZ5D-D+R6I,b=YIU]d5ECX^)O<7FDebW1X5EWV+Fa,<0.cI#T2]2ZCCb5D-(a
RANegKMgO3U=b&aY6eDbC=@@A>#5N]Y&6(P4UWE]F[9<S@#PHOa>bYWeRd[cV<SM
M4GI\c\C8.<4MC@Z=,J=^M)d5#ga7(IC_546A76cW^4bJYZOgea.,?\I2LeYQLR5
(gc>afb,ACNV,gUKe-0;OMZB=:[U384RQ-:/X-7?@QeEf0Ha[VfE#H9U4IAUI;d5
@?+I2f9)MT=eDEZG+04,a9):@f+2=5S505ce@;VL19TGfW@fCH>b:bB6:U)<N-d3
UAK>7cKH-)0d:,f_WQX)B28F;&&+[gQEB.\=U0\aW4>N&B88;d]e;7?[6\N,I@,P
M>29KOVFY#EUF&N)gY5Nf3_f90#/=,4fK?3)&_e-4=9S0CFK=TO1)O^&+TO@1P7X
.8c:YHN/LOTOg8M9MPD.1S,^QI3HXE]Q@[/aU8<(W,TT4_C#HVbe:,A#[J_/.\Ua
W;GM44K.0Z.W-I6>cL62T:US\ACI[C\F7^7&?33E^KZK/5:T)[>YePYLZ//>TBH]
VO:6\b@gMe#C0SN?D#0g(1KY(5FAT[86PCM01W.(Q/C8K=+C2;-\abG:bYE:XF0[
#\cNK7-+XD]9-[eN97_K,P7YX\AVRJ/->I_)--N3VEV2Q?4dBd@D_OS9I<-+d(.<
e>>g5BH/=\Z9OB/0Z2DPV,(Q-0)B&R:=8WN-8Q,SZZS4^J&UfIe+Q6=R81[2Z7RQ
R^SS\b;=6QDLD0+gb-4QKY?^K8GZK0Q78ZHAB5]4Z0:eegaU/+JUN.3+b,7+cHID
Z?7D)#cA>+G;37I<fHZ_ZVWD78KZ8Hf^JL]5V2HM4A7,=9#79P_J9+5POV+Y]P>&
2^=HPWO.8[.F\L@8;;\HP4#FYN.(].C[\7;]-fQf0H[.4ZOa,W3R?>b2=Rc2H2SN
,&=P=e=bG^e1^4cKGCKI)BSO;=9cYBYE2cQ1_H7XZe8F_,=gP+BGNR[gQ:=f0E24
D;&Oa.d7>H_O+JQ=?A#0gLE?[5TEC0OD#T18IA61CF2.:DZ)\-gG/BVK<,LMG?2g
_]UO57[HBZ^4@S[L6ZLE;:ET#IIHDG]Eg,fDSUA4O#)M-6H^,#P&GN(67^C6)E<g
P_U.WdRYN&)Cf74_J7ed@#MQAY1<5/C4F<CIbVQ#)Ug:&:B(Q)2WPbFc.f.SXa3f
M3G?g3&Y>II4,5[UdOf0QF[RP;KIP,,Z3Z[UbP:PD/C4)776(:c.)a.W/_AG-Y;7
a31BULYSDa1a>H&cLXJOdaB@?,QdY._0,OdAdfWL&Q(5D;JFU[3=U,R-I@a_JD9E
PM(;W+=6JPP_^W?]327).Y1E5X^(b6<FPJMA^[EXC&gf#2U0aG;>)+E<]9EHBN[L
[cTWC<WA<T)6\a:]OCQW,7#4SG<BO1\V)(&GNSQZ93.@&IMXHW#.Y(Q;YDgf6#d-
3gHP=Q@4d9f[<XWd;<YN8PO]T=e/F(S\2Qa^S2BH5&STW+V9\K:F317LVQV:be)Z
D:bb\-YSe;LeH87YGS/97P\VFB)60U@aDK@(<-2:VFW)RY=fBZOZ?&1YBAOXgU0g
Zc#IgHKF43BCYLN&e_@7J.WIK=F0G&#Z@Y\dP-EMPZcCD4#GPe.PW#M,,[L68\27
HMbA70AVOKKV)e:R:8eV4^N=&-2#]P78=\03NBAP:(#Z>80<AMK+R0@VQ4G]U@SF
VSN:Vga5#CM:ZdaDca;I<+.5-Da0W6NR+A^>cJC=:))](,-?a@0Tg<b#X946bRb#
W^-JR@LM\IT#a/5]\DZ_aAO/>DN-bXd1_\7\75)KeLJ]+MZ3([=GQeg@BcAdP4;O
WDE>OPC&FTP8CGFB#Z&]YNGZLC[I][cV,D0Y=9XGBLfgM.(9A+S8C1T1\38MOQ6N
?GY[-,Q0[;f7T4EUF-?>aTO]c751O=(AEVDUE)38ZI8#W@?F-TYPM-MKcUA>^K\,
ba,bC<<>3VG]bR_-W0R:NOU8SeBcBZWIF-a1=A^5D_Z68aNa.<_-1\WGOY;_BLBb
d9=Y)G0Ke485Nbc@097a?;O;#[dW_Y18,Y8R3CDMFN]b);g8^Sc@P0+9SXFf8F:V
I=d<5TGN2]MRXQ)M_KXW\G<>[)0(gB\2?4K0NAYe#:dTQd)D\MCf\UD<UG)feg])
1#44G_-=MGaR61.A4)6T;6X6=#X=?]>ee3NDZV1R05B3A)S&G(9Y3NMb2cXAEGPA
f1Q0A,,^;fEAX^G163f#(?caW)c1)8T=Z09;KZ>1[OS0Y.7.^7Z=UP;1WRQSWW?D
-0-GZJNZD?0R2H0(V.RO.+>5a@\DGR)[O@UTW?-[2c?C/EO2DcQVCTGeFT4(Ob\B
P/&cU]U?9RU2XK;bX,^OEP39U]Q###N8#(64b+I_,eDRO=TeJB75=,#R?2&T-66/
TQfJfGI46AJH+2^eI2T\9/[@^O^DU2(8U(IDFfg>=;I0+=+)D&bGYBQ8T_&YVPd7
(DX1;PCZ3F&EWa]]O3c9C;X^,\+AHBL+&HC-aCV@TT.G<LM\RS.#_KO53a).11V\
cdd5GM/<#@&N@IK55\YKH]8^YXdF5P-YK@a&;69\)H0YXYY@-T52bWJ2<[T<WaL2
>Td?2S3]HT>:ESa4Ma/R7)D:E?TfT2:79>)7?\88E_E=0DbObV1-?f4<3g#gSRR5
A#@)BH)B00HFP@G(_3?a2]5gYKJR?,c2R)M7.I?6I,C@Z?417>O(:6VX_?&(&,B=
QXc\4;&XB?F;.?@@M_RE(J?2a-T0\.PE3HO/O\9^N,7B[f]K?C;gGVS4OYc13@KB
6A\@C>2f(Z;+<M>(3<=#G:(^QS34373:_9LJ>M?]SC-U9A(L15GaD-IB7^4,X>UR
;5._S[+C+]OJ[U?R.?C#g+N4C&Y#eK1BGJ9f40B<D;U<OLY9,^@J/_2)A,C9HRS(
)DX/IJb[ZC.V=HaC]@22fX@,Q^Gc]7Y(PH/2Ig3:WLdVd2MA_2M>@3OHG/@d2X_=
ag<DTFOc?bK+>?4cS8]W8?&](Sg(7d6gLVGF>2,ae5?1)[eW4PSZZ^DMNG[Vgg4e
:cJc:U>Oa#,_TMG_gLHa?Z\;<5KO=UXT?KQ,.b>\BGc)I<H;UDM6cUAPEGE:)>SL
RIe(B,&MP=E/BRJA\_GC3beN/:]Sd/UR;FNERJ2CSDI&67LAfRTB1O@S;<99N#d_
2<J,FWCO5+H3;:135MA]dUH4LA5+Q3Gg(bDN?-.P3bN>2/8SI]&MT3[XM&SJ:_UE
L<K/d;Ade/31WAR(E/Z,b]<LaR]bMIHF:DdD-?fOY@@MUT./gK&0X31DVdadF;aP
OO_1REaUEOKS&BU/-PVK93WSU1H8AU>=)^c5K)?;/)ABdOS80cG<+5&J,NYTAO4_
0BC9/.dPLGZ.J><Md(]?@:RPAY.@@9K<Q9&,JGF#d\d[O8\6QUKAcA9e?fN/UMOQ
gDJe/ZTVF8EU]?T&P)WO.)R80#/NPZJ.Q8I6B-?QgN(8BAbG[XdCCf3[SPRb6=O-
^9[E[ZB#75fA0&P+GM_:2bf38UE@g@QeJP[6=1/1I?=,X\[.PK-&8ga(DcUW#^R4
0^f:G@&##T4/27e(R]U[0P,^PDA,_I;d4DeN>MM/5ML&3/:V:)Q+4\6ER.^;XIfY
CB5LJ_b#3^KT9IB2]WP9V0T-]Z+:1B8F#&NeHOMM3Q)KgIBeZ?#D#3T2SS+1f[=J
AGJe+>N,e?E;N_2^0[[]AJ3fTc^T4g@9KU<H\aMVG8PFKI0O9PA&f_.7GcCR]2bA
3N/Q_5<1e^@4>Q^CI0fX)17Q?E&A2&B;ZRcWHR/gcUM#EIM=4CD8?4E)Fa3.S#:4
Y-EGUa^A7#dbOF.-(e_MV];/Z17G;f_[9,AeNW/]36)[^<Q;E;eS9^BYONQ)T.=F
C\dQE#MU(9-P<><B#/KK8&E&5018.=P:U3)/6&7RN9=XG#O0]VKc&#:_]N3M@H4I
BWP<=^g-e/ZI_^(#gU[SO:HOZEd5+GAKb)UISGa.[:7/8U2:dXB\JcN:6I@8b>ZQ
)0J]YI_V.AI52gLW-1)YaZ-@9Q?PD5NCVN1[GECPCDb[;;0V=&HE8E<D78,K,WSP
H5P_eb+KGfW(fa3/c]&Vc6-?MeEE]GcOK[KfHZAgPdG+RC+VICH9gDc\;K<f2K=,
eB<e(\4MLXO_@/2W5Cc.K0_Vf70,+RDO@5)+;YE5Z;9,:98g&>2<BW,ZbfLS,Q-K
0R4X#G64X]]Qc,/=B[2c7N,P)(:e>I[O/R+@NfV;D8);?S\YA1-X<.5TF?SgL85^
K@GKfUW3[D\QeP>d)AJ4JZR[?&0?9a]If9L6W5A,(_CHR8Qc(1MZ6(VCDJX+ZE51
T>X9g9Z5E#HX_:ff)70A^b7bZ9C,(=(PNR/CW3N5Y&#Bf.Q[;60&,Ic,TC4)4)(]
E[>9XU<5X97?JAefVDIV4@1\SP(_UJDP[LDg546,=JIAY+G)2f#&USS8.(F0WT30
8=>g4^L1d5HF>RG(:We_LB,f<##XJg?J-,6J+<;E[R9Q91[^B7a))cMMb;1A4;F&
Q,ZV6KU@@aH_I:aY5#_7R3,@ZceVQ;dZgRd)J@\O_E-/3bT3gK;.8cNL0P9):64,
U7dVBOf0BR?42P-A4QHE6XYf@d+<-\YfcM^1D(U\eT7.GU==?MHHg+YKX9g\2OFV
N?L70::1Q/Z+^..2V8\5\H6PDaX^TV#/->O@1Ud<YHZH4P3IdXM@0VG;<Db##K,/
D<BVVEE3,8+UAXdRZ#d4YR3fYfND^WGNeH?ZMKV@Td/PM7fPf5#eX:-=d=PBMK//
Ba0YWe4P;dPfN^<8DF2ZDXLY3Y)\J[H-+>NIJVHc@WeDS80dE(WY<GXN<WE:<JZ9
SIE6SgQ^53A/\J2UdJ7VL\O-d(P1H=Z5Lc,/)(QMZM[QARdd#+?[,633J_^GbWGW
FdSaa697S6.P+NW@Q@e>\6QEL6d&I+]f\Y2aEb1(6W_Rc,]LCUDH=<_(])1ebTKW
aTN-4eXbG.\Z:3:<JR8bSXX<8DF)&)=W68R;-,S=Bf2+]Le#CBR0^^)(d(NG(Vda
NWM-6BFTWEccIRRMHQ++A+LgO,Q.-\.GYMJ6b1@d=Q:<=1:GD0]>_S:[ag&VeF?5
UP;O0d]/;TW]-</O0b2A(7L96?AGa>>-G+OD(YVK9Ef5eL7b:++d4P@SDE-/AX3D
S:6ZJ@<6S_(R,bgH6C321:F:P=83=.?IJ8\[.Ef(#=5<3:g@9->W2;975-7,;SW8
5L&<0L;XP5ZTcT\X+I52B.ERMYNT6M30M?^.cOY1#G?QV3/9a&/APH;\:A@)O03O
?bF3FHD_E[fPM@TPc)1W<Ge\V]T0d6(MQWK1Y+Z9H33/05F:))ESegE>>/;CaXVD
YU7MPQ4P\f>FYC137cO35@-4GYIWYC3H35\KPE=@VdQ<GCC-^Uf:Rg/WI+Bg[WM2
WXAPZ^_JX3e/W@>#V&cXPVSg>gQN4I5@0M6G_)PSdKgGDVG&<^aD2Q;V=G87\5K7
Q<YSF36B\P&cHEdLd^HGgGb0CSP,(=+<N8FSO:[0Sc+L)WMB/REbN3)=J4L4R6AR
b/IT5X?L&:@b_\TN)[Y;8b<@5_.7E=7^BA5eV^SV?\A_NRgA-QN/6@)#DIR&5L32
K=Y62X,SLE[FO=<<Q]GWY8e5MF?b0-Y)U;K5ISUD7/K5O67P+L;3DK/;@^fBMd+(
;8,9Xg?Z9ZNS9.]S.:2&+W;]:2\(,bNAK/EXR#dF^:P+SE[g:]ET=JYPEcaWA,,J
^T&@Jf#RKUCGN\15E<B3H,b\KQQ/C?JaEQU;O-RV\0E;4(0KPX(46;4@c/NU]U#M
eQE#JYVQ5a=:^S)4R@.).F#Z5<Q@@O[&ST:gdT>-(bMLG-,D8U.P.eT>R_Z_O:LH
@E6FO+:-S>_T>REL]LH9AH2B\ZAAc;LJ#LfV/3P<EXW0/6L&Fc0>/<OFY+-4=TdF
5,6E)2@D1Q0?6Y7UD=_.&Yb72HZOOJ7F4(:1WRMEb\-=/N4TO-/SV\[#1.fc4fbA
McY:3&UUF5B[A:59?]U9F0FRDD+)E4M\dTM&+75#21PO2[<JPC014IGdM6?MUaQU
=;/EP3F>G)#WDPaG#d9Y[KDLcbU?N?HBQ\=VgeX.)@dY8cZ(@Q;U^OASVQd.2X\e
RS998CP.eG_T1&0+EA],8Pc,)W-#7GgJJcI8H8bN)=?_:ZO-757ASaNR-=W5X\g3
WGaSeO=]g#:O(YPIBZaf2_F<PARDYfa8SX/\;HJ4^beQQIR;=8O:LN,[eKV/4&V2
7(DM<9X49>+NGdIe5]R9TTA5,c53)c-]KcDf1><87^9UE-&[]YffBRY4VZWc34OP
E,FbP#]V_)&CL@K.Ec7DATN#X#e1_cD9&-FX[IJ4+EJ4CB7,,)K<[X64)gU(Q6<g
N08e5ZD87WPUc&^#ebZ(M\VWfM>&=88ZbDaYQ=N[Fa)7^)Y_A.L6(E(O(=)SO_;;
VQUNHd,f+KgM]&5=6Z,K52JE^\0ZAbH;e76#<b_24=;RK8A<:D,ECO@2ZCO]8-Ne
gb\3FFOW_3I2J.;@:-A7Nd;W2X</ZS44E7ZcEd(=:+;8\<99GAF<].<gHb\.YWOF
Q\b\=2\1=U179<O>;4&@MfRGfU4de0@VCR[C2&\F#=^Ba\Y&2IO8f+4?C2,@]>;C
1DR4,4B)@#T2ZY2S/Z76MT#6)Pa8bOT=>AC[@)]B)c>fcIQ;,aEKC[0J)9>\^0+R
5S86.H+#)<[LO((d4H->O8<+?K/=UQ_caa?E6[T#3D,S(6[E=;(Z#5+D3I_bYVNe
1A_F2(INB<.NCOR<@7,I4[N2HWG230VO2,IS>BO-T/FH46)NEMBLH[&6EGLOJU.5
dU7GQI&Kff?UE;5<S,^_^MBD&B8YBF1A,[P:Ug]J@4/B#SJH:WNRN#GDAFTg)+,Y
<30,B]:,dTNDYB[4[G/[6#)gZH]7+[O13R8C5WA>C<e06]E(Y<EeGZ=bgeQG@AZX
FgcDF(X2WBPZ?2J51a#fUFZSY)97>K[DK=Gd>[LB.fNcf054gaH@dT0(eY9G6@e&
VFgD@8IZ8,S.SG-(G]aBI&45.65SZ-<@L^EYa@Z1B9BRa?=d2DaFM?K^;#CR4?J>
&)c#=J]g4X&J?(XKJc[+?HKT+L4V3C0ZA()>UT)>KIU\/O5;\NOeS,<K.4dc4&D_
-TPgW<<T(6&eBW18aL9=-#HcS_61]+9IJ0#e,ddD:Y@#XTE=8KYB8O>JBO4^P0Zd
3#2U^H<<Hgd@<7>P/a5C\NEBK8HCEDC)>\5)bHEAR_[=63f5Y#?X9K9N4HXN/Y5#
W?.P9<EgD2U;[^HAUSE-5OO<+O)7K;2&6BN22D)TNX686f=R/.0HBZG&@>^:WGZJ
FH\TTGSb;UT=ZTFL.f<G>44.MS<@UI4SFeF&F3^?BX)e8KM:Z2XR=YDNUNE69EDO
Ic^NccM^dEa)7FNVCK.4NcPWXN@5&]<2g,VWbKf05M0,UNcOZ\b3UWPW.+b6OD-2
e\63(gHdd\QUGM_..<eR?@Q#OG9XK<X57C_HZ.aF,CQJ8084Q&L1LcY,EGgL,TJa
&98J.LTX2^c4^:9:4IXY,8&CL/I9DJ_?dEW?]M];Y.KbM6[Y.5:>:NfC6IS,c<[2
0d6.[R9J\L7<TE,8Y/(@]2Rc5B_HA_]1&1Z(fHMUP3B?&[:JE@]_B@M_OgR:3H2L
LJMcH\Fg-8_e<,Q^F[63D_UV^1<=caJS63@^NA)b@7gSD,&bZg:U_ff)Qf<D1RW1
W_a<^;C,R3Q5Y>cZ4=SZ+G-&_/e.ZI)g[7&[_69<+CD7;&0_B=4<c2GU+.E3/b@@
^HT,9>^;)77VN3\=a/eU_b77\f>(4:<:4+GAIFO,68B[fg(-/^AKN28C=[S#PV3e
TEPg/J[1b3]2Z?;+4/dU&dQ<FB>/XL734J9f^FK5JNagCBOB#YRIGZ2T8<[)^_,]
#YVFfeMME:ZP)RRV;3#^9E@.D38+?NRRYC/YB]LaR:QTIf;O1f..bLYYgWK2U=9>
DLXYdV(T@/:B&9=QaDPc(-11WU0/gD.OR.Z0\L8Ua&,1>+T7)2>/^([=Z^Fe6A?1
WM68B8TF0\./-?8baTN9PTX2^4L.OFLKEb2+H-938,F:?@]Z:B8e75I>UI7[]WgK
ASU9(++8P[T9bCDE@S=Sd2aR3a]5>?0@FT+bM\@2LMA\bUa<X8^E6MbV#0IV)R9N
;G5CZZEd_-V6N(08S@9DgLGb;e1&\gOV^Ce@26\^?4^:I3J.M066(-#,M1&_c,;]
b+bCV:Y_X[0W,aK\deA7dW38-,&:/Yd=<#Uf<-6O3405WgQAHeA8S>41P=[(DC=U
M#12Be#agc];BXX9g7]\g-5NV<TGJVcJCc&;U^g,EM^&aQ9fB;8S?OF[d0/g]_1G
V?INMUEKQ1ICL=9HA/b;VO4FTP)\<P^:&ZNGT9f/_V3R#2^N&P?RW5b^=b_O0&&;
@HA7O0RK+B\11cF9N92e3gLMB;.f\8fE:1f&XP<\^KNW(gE>X4ZJV+S+B0<W;?gG
^?PT/F49TT:.R548,?TV9#ZSG/GF)TEeF#PM906E,dOZ0K[+HY^7fKPH7b(1deWE
]4OdXZ/]CHVU^IJW4=+ecB-KNA7eU^^]Pg5C3ZDYRg9E[LaU^1?NV&0>G.8UH^<b
4a\/SOZ9?[1>&^_VLPA_aDg7dbJOaHB<EUa#<[0:WSF/)R4;[@N]Jg>N8D#V36CH
:U^,edU=DK0[E<^647YbI)=G#>_&?Y:C/;8.2a039fd5dT)JIf<./#QV.eJ5M;QS
?UB.EQ:L[I28#/IZd<G#+=7V<R#/bX.N4ZK9N9;;WB4BS\c6Q8Wd^Lc50AA[DY3C
d3,QC&,7OXJ]XUg@UEY=[\K:3T>D[PZIb8b=3aAcSKV0Q02NN)1<IF(1b[]18JI3
b]Y-7?)M&E[R#ZT#/71YcN6e=d,Ta[M7(Z.&]8C)0MD\7RN[d#@_NZ)LUCWfK2VI
OVB8Q;IQN?,1VdJZ1PVQfSc@1)+=7aWDF/V/e3FDT^6PI,dR3\[F/.SRY(D3:-P4
]#W+@g+;C1#N=e/K3QC=UM[\B_S-YM;]R)R1=>3#]=PIJgd=eMX]>&>QB2E1KONc
3W\7@B)e_8b=>V<PI5_JeH#c0I_G_G@Z.U+8A&_Hc(W[PZKU84c.VK8?96@_a00R
G83CN(,@:>)J7XZb?N\g>5?4GFTIK@<3D4HAX(_-9cY[02[YWdBVSKcFBW?4.Q<M
^:.HCT2>_FU.8[M/fH:KF7fR_Y>gI#U2]A^?NXRIK^NLXZA^1;6IPCHMP6Id];,S
+a2-#3TN/.9B[9gQadYU12Ka&^a,?>d?_XH3ZEBTddPJ1>(CAO7F\@+c;0NVK(FK
WE7/Kd#<ZE\WJO[&S3=U7V(@TLN.JG(N+5a>;&-:Fe4A]H>ac^OZ]&ARCTPAe)1F
aJ:<1,&WSZ0&#Q-IE7C7UAU0:DPMYZPc7,:cZTMVdc[R?GAO2@<,gQ27E9?9Q0?2
aU_MWWHIT:EabFW>[1:VVU:R#.5b@B4MZ+]_>V<,W.Nb@^d-)7S[3<8-aYD2,6:_
QVVR&Ia#-Z:fTF4GC.WbXf]66+C&bX=QW6QQ8T;?XXL_PUJYb&8LIVUGV?2[3=FV
)S]ST@M#L[?d-\a[5F#,U87?L[R>B68@J4=XgRdg0<QPDIQ2^?I6+,R4d7,[PLe,
DK1J2fM29&&aIY4^FfY7PL?R0K@E.#aK@N/3P]-QS.12L>)VZH5<CE@Aa/2aTeDX
?>7];&_cL&HNSEE;1&\1>,\eQ-0/g]753ZGZScg_?^dUM]&/M3QH<daFR?=PX)26
,TNb^gUd]GRJZ9EGe>b4+g4/WV?9H/C9:2164^g4)\U2Z9L8Wg]F08XA#2_(FSHd
3ZaX:VA(VHbNMU\0(SB[-?7Q134YcLI#0Q/O\fN>@\?Tdc&PE@O]PZ9B)>40GLQ,
:)R7.^O@LC4PO&D?S:Fb(CX2)<5U2OW;[=S:KMFAS;5FU^1QYUc/M?U#FF?_9L7E
a(L-@ETa,4HI?^c6.DQ5<LHS:_YD-(gFL^#0SF#YCRR,.57bL8HA95^a/K/d2BU-
g8-R+XVR984S3;@G;OUXQ.V:b0/S]^5T+]OLO2YXd&I/1)O?G\7gZ_d&_(.-)I;;
Q03IMc@DTde3J_,C9Wg<L>;N@+=(Q[754Jd@9AUIP=ET@/f^(&/PQ22-WVUE9/;4
A55?WQ#7Z)EAQG^bZf\A2[B/ZXJ?-L\8\f.N[YN2)c.ECdK(LAF9T7C9cEaGC8a+
<=)c,S3U46;WaA/\A:^eN+=-9T3K.J/a0Zg+\8.ZgI4+C-fV&D->2gT221HU8UU(
ABRV3\SVN]WBJXJ:e&/FLWa,5DE_&>:;ZMbIg.5UEcf[:=8#76P1NK?H8^Q&f=Ie
^ZP5Aa/e()0V/bNI6]3QWS/3FS?^gV2:OW/=Y&d)G9<(-]eD[2bcSX\NCbM,62GE
.3A,WTBNZZ:/TV3@EIFLZSGFQN18&f(LA+O_SH7a=[.a?U+LE[Z?6c_Z=M7c-)8H
gL.7V1^<5_76(0VE62Y<(1OeEW8dMUI4L18RaDL^#=E[ODZcKGbSXSaIVbdPX8#Z
L+#gZ8_/PKJ@C#<1#[/G^OI;OL(=QU6.J,KG<.\>B9J=SBSOg#d:F?Q1L1:0BTV_
A,4QdK(FFQHU<)KH+L;5]d&I(-KTC5?c&cK#ZNP21+BK3TN<?)3c/MK5N84fUM[>
bDK3gQH,OdKQFS7&F<IcbdT7(G0PEa+aF(aIC(#Q,7b_V2(ffCKBX.6-#GCH8Y92
DAaTF4/C1EHJ9Q9,eHNd^Ga_NR&X..5e]ZXWV.&deK_S_\d/0g1G3P.?g(ZWcKM#
+0LG5<6Y[4M5]?5NT_DW-9O:AF6_gR3a)1P.8NDWAY?4SB&5L;U?I[WWgY^7N[:a
Z>9=/4;7H.7HQ]5b:_c+,V4d@GN,^TN+\]3CJGS[6Z4?cC/RE(B<7JPOI\.@@CBO
e,B8:._JVB1?+3<KQgeS_5=c@bK..4bQYdVZ+<N.D<,bZLOE,Q+aSU,WGY@^MJG2
g[9_6,KAE2>)&Vg?/CC-fO)B3.RVeVR6/NTE/0>(d=AeNV==AT,XQY/XM7LKUU?T
.?;0<-fS9],YGZ\):3(@^?/NcU6A.\YT2/TDG>]4/>Q&_;.Q@V@>9Z?9fbKP50.=
8dAf/-RdNOT@?>7R3+LR<a/7c7BZII6@N2(DXM3gODEe:(QJXZQ?-&)aRM.BLYf\
g#SM83VI=b:WgCS9b-]1_=]@Kfa@6CPKe@7f)[d;->DI3F6<6fIN:DVVU2J.OIYT
193;<daeQ[ZA?YZS/dXIQ&CVU=^?][#[<UI047K18EN,C,K:+Q978JS4G_eY>;81
OE&PI[G4U:G;/BU@D9YT7@E-\QPcSSG]LBO:/S/F\JIL.b:Qb&;CM_Hd;ICIC#Ya
Ce]<.1L[)PYE5[B>WI.4TZN_@3XOU7^f+7YWMdS_5fVa3V8ZYaLSQ;7)Rd;DX+\b
)H@LYYbR^/SN91\#b4Sef).-KW:&=XbT[+U7a?C2fX6Y&NPb/Gg?W534AT&[Td@R
:KT1GSHPd)fWWYFCPO=T@J[f8aZ>afO@8>dKKA1(?gGe@Z1;9=TPePE2AEHaVMeK
[Z]2(I)3@_cE<Y82gJE;F.9;9-B7G(Y(.HY5JdFDbQ:8#RCUH2dLbFZ,]PW]c\gK
4D#DGJ.eF:^e\+)eRZK3P<@+<Rdg^\1B>_KgHHWS:HDXM4ZJ).4_L(I\[4e_WU2(
@PS@.gH5H+IIEg_J@S</ATEeQHbW.@A.+^<FP>bZZR5e#1,]G4gf-5RPNMTL]K#S
O#=fMb<=+)?]^RM_RdEY2G=?.61U#5#&@#/_990:_dfJ_52LSdH>;V5PTC;;6;6\
(Y3>IB.)?d=gbgbIDgc+]K;YVaOB[Pa1;8#aeR9L1a?J@T38+]_/NcY_6&_V>OfA
7W>^>19C94g;-<_KC+_:_M-9[-]P6;N?79:;g.1@967V1bA^7Y&OJ,+7OIZ<B@E4
W3^(B4cW7E8:D,;34)a7G)M_[_]<=GVUbW.&]?AH)VGTMR(F1/QU0(c#HKW_6<N\
_L=DBC@3a5aG\/e/:X1-gKN#\CNP8O_(5(WQFXW&7U;9X@8P79)_>23GR8.L.e+<
6gI1Q_J7Ca(PV0#U\VVR_BH3bC/,#F;TM[7+GG:;;QfIRJ.)2MCb7e4;b:eKA,EG
d[HPL>Y2(J==I^8LVN^fb[c;1E+.Da>5,/XY[A0Hce-cO5dWGW>gbZGd^L@0/AfW
f;AL:THbd[\ec3a([F@.FV)J;D](88Da;@C5+^R/g@[WYLTZOAUK2PR,#NDQT44[
]9Z>7(VeII)3+U?.WbdAFbfSV,FQ-YVR:F/Rc])+I3)a8KN-<B72IV_&[K>[1PQW
]+F56=W#+TY_,;WYSQ3IZ7)?9\V)HPG?G3YcH@3cf1)[O]bE2U^R-#IZ/W;S<4?Q
&]Fc>T(0O;)H=-_:5IOdXI]8&270SFP96g>g/]>24_>fN_aZ5VD0Wc_0V7:0/SUC
\EA[K8cAZ;)<@>A3RgASRGVNXgA^b;3^)a&5A+P\=5@KI+gL=gWCPPe5fIUL##_9
eTXS\a[EXLQNG(V8AEF<Y?>]M;:Z]JXDB&S,f^c^+c+1ZP>G7(32f0U5<?(:YbA,
/.XK6;.2<6F2Ia&8ZG9;-Ae7e:>V2OJD^_;W<eL9[V<TXgFRNO1WKN=6^d&c[QIg
@J_efTeZ^0T:fAS)6(ZH@NINI6?PUCQ+Fea[HXYE>fI87HL&f^M&4;4R@bF+_.Of
P0#Oa><L(\cY7[QARcA@33I5[4L4&V=^;G]8UYR2ZSMI&HHAIIbF30P@fAOQ\>@:
N9fLYX4[+I#]e9;BYSRQ+CJ34H0CM.a0/d#9KZ9>[bZTF/@O@K(VVFQ?E#7,O.DT
Wec]&?SHdNP>1OE@4&-g&KZE5g(6?6/P65@cF&IM.B21Oe[M&&6?^\-\/AE;]4DI
@51-QIK/7C\^(U6cY0HgYT](#Nd&fM_,@-e)IDV=+43^GB^1AXZOL7EU3NRUg1-a
)L>BgMKV4aY:K&^VfF:0J5.@IF2^fL6a>c&PTQ_F[HQL6da=0+I]GAL3Y^;O5S@8
;_MecIbK]&TFVd#]@\@Td8K))W:^edH10c+7HVDC;U0gGc+Z6?e7DX1fN1].&I]>
+J-H0L?_\KL+)KTGSdL[8_32Z+OeW67(&3eSFSZTgY6M13-4C3?K)-M4Y+T.TF>;
?]:RQ?I[(VeE>KX5[=_dLA,c;@2a<BeCC5+#?c]MIdbg5_+Y2TN:@^dA094DY8&H
)6NE::>0AZ430C0&gL^D+\.J:9JOgCeVR<W0R#c#gC-=<cJ,YQ&;0EICK9c+-FXf
(_Y1T29#.>cREW-eX]9YUb@3&X4.&N42afU/YCGd6Uf)UBJ:7@Y_D:F<)[gRcT@L
VeA.;dKdb1G.#1-2V9Ha0F_S,M;=A;2)&19a82d4#[K71fZBE)f^MCa4:;MR3T-3
#PeGZCWcL[L+SeW1/)0BP-BW\eX(?D.=UQ+UF:#:,bA_-XFD,3\K@>]U;-g>2B>C
D@CBg?8,P.X5PCH)R,&:5H^\\5b#/:K.I=0FJf&CXOJ\JIb4)-6XQA,>2X>Q8EWV
\Z0VX,bLe=7T^J(UOTWSYLO/aJAN.Kc0ANP0?II9_?bg#RB6PA,)<f(LG[e^4&W,
DV.RS?K<>UA3Gf8#L4e3(XTJ0Q2G[:5Jd/Q4MEZ\JZWe+UF9f@;2OT\YXBLFAR6#
@B;KK3,GBIS1[(O>](MGU.8?c/YF7=Q4;[0(DBXS3]FE4(0&Sg7+9;8Nf8Jf>E[A
7/9-L(O8Aa]6L\=B5J<^GKOeS-1TW-MgGKRfCNWU1EL[8eTOK:-_L>R:<a]1OaN\
43GKM@AfZ(3E.GF38<T7_@8f8,cRdQDZf/&H[+6NE0d&P=1KJgL>UJ5:M^#cCd8^
R)2&RR-B#;ZWBFJFZe[7JP_Ma02#YU9QB&B.[5/LH:_VcdM,1&/_->IGX,Xb,IWS
?AEVYd_Z^7CBJA[FA38g^f4c?0Y<7<_&;G>K.f/_VfS[&.TSGGSD-Kd7@JCWb/^A
DNL6LP-b_/(Q5P?XHQTD1AKU5SEH?-#=1R9-/?SB71ARH?(<_65]>EUY(?K1XW3\
K_R8-;WIM+EEDA;Z6Ge+agfL[T9:X>_O.?dfD<Ye4S)P;6>ZDRbLW9D9\R-SBU[0
AD\I)1Q6,_PJ?I]MP2<2>\fYQTc<K9;-.B_SN/X]7c;d_2J4f\N-[G?X6QW;UD,)
L2(R]VY\,4KAPRe1Sfe;ae1N.K+=ULTO[RObdUa@0IHN--51FSDF6??)f,5.bA^V
_M87&)Ac8F8-g.MXW.5#]\,:/C[A3B\H(3dBSJO3c1/)aP,UPN>PY-H2HJBY=B=6
S5HO_WQ1&+MW;)MUJ]>bM9#B\JO5G#EcS^6c4+L=fD8(YJSI1\52b2)H[#c=2@N&
URC-,d9I+:cdT8P8>fR/B6;HT5V=5a0LJ3SIg7QG(ga<DL9M??cd6)a,OZYF84Ce
0\R_4Ba_MI(-V],0K&UU^R9G_?,QL&<#=_3QS])^EIEgY?@C&Y>I=&I9R=c+1T(I
7NYFbS=J0WX0Z6[6=-9\:c67XSgS?2MH@GRa1@<7R]WD][bK8+DZ3]OH;0HMY6]g
V(L,]]d,,T.Y&NEd./.dOb<N;LWV,Hg&#G(F>f[-4CG6_Z,/AK7>J+CP:PE9.b2c
dIIZG2BQK;EGC@-b6L#bUV95Rf3UL8C(EBM<:M.=,b\L(<f&7dI<GGdW)DTe?<ag
RRZQX7XQGLQca(=?XPBDV_O4[fd-Ba0dDVKR:Xa)Yb3+Rccc18R=_FD2+:4]UHW9
MYJ8L3G<O0UWF:L=H;e78/GeT9Q?S-R7ISRV9<W,L^S#_L/6:cKWFDg3R\c^P&;)
2dYOaV+3dbXN[[72P<VX50BQTA@g])c&67cB^b():D?=TH.N@LDTBfDK19C[QP-S
;N:bQd\JEM=?(6/^0^[8MD3]Z;#;f+a]eP4RPPR<G?A\=7.Y=@W92c?A/TB<4NOO
&ZfJf-VY>U[PBR^#OG)\O.37g9JC=Zdg-=7^D-.f/XQ\4#ebDg&ILY>/NbH-ec7g
B:G04#XdXG=&Y<E@=5ZaHU_,B,@dPS5R;Q_3]XJ5BL\cagR9)907BQMZ5e6NDHLS
0F6WI1+DOV)Q2#5WL+E<g15E+bF9eNC11#cAJEBfC,845X^>371MfYVDcY7.Q(1>
;=K^cQI1O?P\A1;VII#?\(Z?4Ua]<RDC]e>(/F+R&.A+46[))EB^8/W7R0OM/G&T
cRFDW)R)P9=(61LKJTcU1KcD3,E#6YXE4TfB[G+\Q/1-XQb9+HVNOL3:FK8<LV_)
d?g-(#OR;:4Ge+(C;O(DU1g:Sf[D]1OBR-V_GW?[9R8;Z#X];MZ^6W3ZOVR0(X?b
dW(+C3/Q=LM\6MNVcdSD_\H@95L^_g:W=K8)1FP]E4AEbLV_UcTYF]G=)-1=CP-N
QNBP<^XRZ:F20dg#EHBO7d_PXRf\6+4]a^>&EI21XH.U6NMNRP@^;EWaB<9aP+6e
2?1TF(YaOE.(@R5SZ/DSAY?,R(G?#a&^W+?_0]EO4LPW.WdbVDX+N\3RGSXCd.cB
b8VI<LP.3e3XAb)Ycg#<d-TE4+W6Y&FHB([[U\N2M)69/W)D];M8RG/JegE&[Q?T
;-K^]Wa.,C[.W86,7de)]D:gOgTXVI62:A0FOeHJ_\.W=F:>KXK15BQBS^AK-@_b
&V^O6_>abc]SG))d3Pa#O8?QJf6A3G7(a:OYB1I)d.+<WdfaS]FK954-cHNU]U7F
/]5IU/TQ\/bVV5ZKBE,PeI+gODL@++0&-RTGW;<&6I1FYI@Zge]JceKS9P&:0b\L
CG-2HK8,RBcPd+UC##4a46EP^?,f3L?33?2bcVH;4gAI2eV]dC>(@7S?4KB?6g+0
MDJA/Af2RF;WAF?[Z&c3VdGDD-NeU]M1MQ_A+@fHML/cH2_WMWb5d<5(&W-(AUQ2
cbY+VGa;#Q9UR?,U([&WfE@^MQM89#K=\D609cVe[FSE&dKWcc^_J?AX@7UM9F20
_#Je>,/A];?eVHDAS?7L\JXC.6gYFN8L4/,LV<g@F).W7]a5HdRBUF:OEID0:\D9
],c<TSbQ50P_Ub\DH8]&RC7L=4.QZTGW64\)PJO4aaB1D<+beZ60D&&O9,1N+Ncb
NU5]1X(b@C:KG(Ta=F.<PWJf08=-O3,=3N78+@[HE=N]4<M:RG=DM<=fS_I5AQ[g
-JGZJF,[C2F6CV#==M^:<6:#@D:=J2eH0c6YGH=^J]B>)a5?4=Z679#:dUb1&\4[
QaMO2D4#Q-d#N&;9<-RM&W,E+O;+<>Q-)?:R(]12]>L1O@X&U>Y?dFaU_39DgBWO
f=\e_)?b#EEAMRf+TN]2Ua6YQNCN,/VUdVa[e+,ZE5A5CL6HR.Y_>ZE4Fg:S9C=I
aO48AN_,Jc1#2U0W8RIFeI2(>P]\34c&\A25+N<bJgC^VH=@8,RT\^@D6;Jf-5Kf
MF(ZKWT\I_e]4/?:EB07QW-bVT6gCafe;IDZ&=ZUMVCHQS[&EEB^D/Uc_<;?)7B1
SDOFOM<HF>H>OWI06ad-R5L[b],FF^[CZG[;OR,?E)8QXL#-4P,S>+_PDg-S6;Y.
N,T&0?#XYd8^8eI^K^AKQD_8aTGPZcX]d&@Z;db\DdA;75N&0;,]_RdT8Xc;KMPD
ag,^Jd?:0O20>]8/80.9GE4M@ad[G8CXM(+0_;eC2g(3Vfd-[-C2fUHFUD,D^3S0
@3c7(2_91Ib\bGb6&IO(RCfERMdPF7g8T+=^7aO\839dga,]N8T2=B86N9(<7:14
;<R,eOHAVS-B_aKOPYa;U>gL)Vc5EA1.CBI]-c7?]EF_6QI;QO9&6#5CERN2I4A6
+1b/M?.-(fW(?6A>Tg]URC>bJY?SYFeU7VKCO(2Q2B;;Z+H]+ZKD/A0aH_XAYd>d
+f,YR/ZWSVa]-^R?.f(?(.M^A2I8_7>J)37G-@J_06H7IXf;G/R(IFH^L?/LJ9NJ
-(IB>e0#LD0;.D(LBD=:7Ff\YR/9\:M2\JGYREDI7MbAWTU_>XK16ZO8VHeE>+aC
:IM0bbT64===X^;8N13J8B0:RQTKUDCd#?7X1H?NbO_.cQ#/\HV=[W<YFV;;9HQI
_N(#YIIYU-88<bg)]F:JN@]b&RP_P_b0P.Og;CgU4/;eEe,_-<ZZf0-G[9>EQ0g^
=(18V;0C7Y\CSWA[;,-^L1]#afGJB36JC+=E)eaF4Q524.Y1?JcRZ-)(\^OR0;DE
84g@/e<a=5:&)X#g0b@GBDC;SLCB+OT89(+(GIPCOU9-=H,)QFQWDUPA/.g3)_dA
W#51ABdFAH3-gW04B7DX_9T<O-W-@/3D^dCE[JF\Ja_=P\84QE4[J=P;Y8a[_+)O
(eO6^P0^F=_QDEg4==BQRV_8C:X00S1+KAX,a?bfO98\L_gVgP3+M8;JMJ&6UgS=
1;Cg-]ITU(g@JY^OCQ3VTX)K?ZQMT7H&=)ZQ92I\^^G<R41SY7H=9=AWN(C,#0Zg
7?]ME+0K)/FfG:8_;NU4)+Y-_6CSO<B)5aWU?]N,FA;<&S,10&^,OGQID2P)V-?f
g4]GWN<FRa)aHMd@I9(^J2(@?]VP1DY+dDVDO.e9@P>/b=JLXad(F^fKF-6YO0HV
7cY8;+2d@)>NfQEGIU^9J4KGC)S8a^HWHKS1b1#?P]/E?>E>&fQ6aW6,8c.F;ACb
KKBaVUP#TQF^?2X@b0I8C>EC=YUZ=a.=g(IEN:d9NUN>AR#@Z>/&E=Sd_g8[X9;E
U-@(92Q8[(fNbSKRPE8-GLf,;\D/8O,\@@W?0X,NAD1=^_X22\_14[REPF]&3)4c
_.XcD_YcDS6gSd+1K.eXHNL.R9_W+7^=+DRK+e(J<BZX=5>WV)?]b_3B2MeNf0[g
07IKTK(#N[,7&EC(Zd[0F9DBb#4egAdY0,H\VNW@01XYabU?A\JS#I+3YY3<VWeU
4_Ce7&D73XG?F#MQ6V0XcVO:e-.G/2U]>X&?.6<SWG7,2P5.L7Ac-g9g:76A)?17
4^>9,C6eJ<\2C_2@0bOMTUTRSa<eT6/&\5[<gg\,-MD0fP_d<fT):XR)@_R8H4e8
KN@6M,H>b62M[eG1F@QPAVb&M/1gCgD.XV.5fPYBKH;bK#:Ec63e?Kc@9_3.,QV_
XeXRd(OfT17A]Q[0F\QdVCCXND)AN1OWYJ\K6GG@_Ue3+(#6M&/5-TR?1L:H?3(M
=56Ab&7OR#K<28HC0^TM).1,&]9W^0M=&^^KT^Y1fY3c[#-9S=<:9<&d1<Y0@d.=
)_/1&\/0;9X?F&b5ca5U&aa)A-)(3F@IJ5/5,L-/QL0fH26EK_,YU&4;,/;[60cI
^N>ZaO-I;Y1(4e&Y0,T[+_HAF:5g^3H4Nf5##SJEYZ8da?=#eT?36MU;da.9)8C@
8ag534Z5QcD[AS/^LfA2?9DAQ@8J@Z@A787#JeO<-DQ>Sa_WGK>4d;+S9Yb]2_D0
;B-4CBd?2g4W@G>0IRc>H+a=c[c,V/LL4AD,J#TAKZF?#<5RG(e/G8_H+=.MfR44
Y=H1Y)Sc>WNVQaZZ,RKFEV,Ng&3:F<H3DUaPOG(.BCN1V+:6RD1=_TcT\e//2dYG
APZRN.VQ9LdUJP1cW^0<aL5C29<7B4#bNAMd=S:\BY+SBLegG@XI5KZ6<_bP:G0X
BC1L(HW=B@DcM#SG51dDYcA34aPO^/aGWRUKS:_S^DK3+BUf#OdHX@I_Za32WA@a
ac4;\a0&PY7.g_5G5SU6aacf(0c44Ga+SU]AR#;/2\Pf4&O</B/^T]f__03;e&Vb
FY<P6/8O4fRU@#[D[1R(f>7=d9<-E8J=(-7\?75cMJV<=S3I=PTY@\]BAZBg:YT#
b4a8CX6RK3R8>(N+^/R/5[0IHMg9@cRfB\K+M)S1HNb:/,JVC;AA4Jg^99DK/XJT
SBILbKHY=c4V=b5JZ59-HK8&DOV7CE9?GdMJ0^QR69I_03(fD6M=-&J\\de)2Y?5
^&S=A_c>dVbX\ROe/5(3TCR^G))b,MS_@@V_-8(K@3)3K/[7+:4IXMR7Z8#)K>YL
b/?)+S[J5a@f8](KeAA)-PXaCRI3g;3cRN9;eb-SCab(ADEWO:f=\_0;>9-L&ZJ;
7(W.:@1XeUG/W7?.WS#3VYaAUD-33<M3XF=E)7L6/#@d(I]0O6Y&^1)X6L<D7>KV
W8N@_&@Ja3=&dOCdR4R#Hc>AP1N(\MI/8XEeP99271].b7FS\g/Pf(+19@?/SRL>
-.DVgPaTS7Z(MF5D@c&]-&EQD?SBPA:7S0gJGEJC0&fcNJMT@XY<?+/<0.(92#bO
1,<:.D)fcG+U_?2#@V.VJZ#827a?+WW5<COHA+>W2MaEXIZ=7c;5Oe+1BG[Q-gaW
Y5XR-Y:b@)=)[3b(;gSLA6?B2a\L9NA)FXQOD7VI=HY#J#Y/L7LJXcFY,5,IW(9=
R.X-eA@GX;W0^32INdK\V_T+VXAM<a?#OPZSS&WGVK[V_@3VXX[dQTSaID&fCE:I
XVD1WfDPH]E9(B:;H4P&7JS(N644X[+Pcf.8Vaf+Z>fR+^:[4J4V/6.c5T7Kf\W4
e5LX-R5d/6SF&Y5[OK8=_ec&5HF(,R]cG[c;NfcP8)/#IPgB;<U72f<JJP1A7U_4
\H@LBK\3gBQ5.cgB=0g?.X+Td5V5#E:BKG>Kc)\7b]OLB[Y>d;:-:M,]/9abWZDI
W=<I6H;1AUXe@L8YLbWC_WaG<feD92G9@ARYD-OX_Gb:#?8@.+SNN4SId;6b_A5e
F:J?YVf(WVLB@f?./gbL\^?Y=F1<56a,ZfbgJR^AG9GdT;RdN(EBMd(2:WSEa95W
#A?\^5I^<HZeJ:_SZEA]T=&7c8H-4d<VdFeUHHFIQSaA03),-),+F@X>_(2,<R?=
ef+FZR=N#:G1=>UC4\I)-?6@CG]V&&8&4a3H-3VNX^eP&?W+e1G;]L._gOHe_aZ:
W>R>C_?F(bY,@b[&^6\N7W^5Df1Q)O:-#;0Y\7W>UF#4^F_M]FHCS#GbFa5;(e1?
9K;Df)4QLB+UgGASCGK[AB\/M?#&e<YR_PV/M]4^BY3W-g]2dUO^eLdP3?f7fg=f
g1I)6(b+#K.]TPLAUBYS3Y#,XD85[gQ(DXVa4@58K4[cW4UWd7Va=eDV\[JG=J=A
T#PKa)J@7LCS3XROCgCb5,^=dO#ea5B6=F6EVI;@@=ZeMH54U\P\@\WH@fd:I4_2
&#^Eb)DWC[RB9&f2>5;?DGT(MHZ:0FEEP\2d)LR-g@-0<1L,O<D7b+VSJWbV-Jd4
Yab3g5Y/1+,b<N]6[LC-1-gM)HN.>-</NC7=@SWBUS4AU<D,[;_[dcNH.IQ0aA8/
&..?^:Da7]U.V#-[RZ/\=F_Sa_/(;1,,&#3YT+cOGJY7KDQA[[/0fNbCG95GOD+a
d/8/W1R-173K7.REb3O+Yb9fg=MNT>RLSGN,.(P<.IV=M#Va?8]<aI9GQO[f,.VS
2JR.K#+.N>JBH:EMb+#^0E1cbD\M3ES&\3gUVUWbZBC7@XE]=5F;1^,#^dc,d2<W
[B=U5=W/g;,OdC\J9X&_>ZT_e^5FQTP]7WX7fWM4A3-+<X/XNFf2CG3^-+W(/H<c
<+\;G;2S][]IJU7bKW3K7eRb=;5^KRZW8UZ.KHT\<=5&,#d7AM<33_ZMA78Wb1NH
-MHA-Fc:SDRWKX(<;8HCba.6+4KW;((9+e8?76=e-bYcP\]]+0ZPO=g<+XGdL.Ic
]8Z.(,4_@L^([23=H]ZG>BBc&,]<P6=C5^D)WD7>OKXQ=^/[1Mg?a#Q)Wd#Q^LF<
Od(G0?L16-LH/DNRMA3cE)UXaB8PWcFON&-<>U(Y+6c1b\K+2/=d?(0+N2f/-c&c
J:XA4=Xf;C1de)EPS.?<S\NI_eP)10EKd/&FB9d9+H_NS+d?.RAO2>P[:4/b,@51
<3AU;+K?;D341#FJ@QD>X7PeAIS0X9I#F)SEV\R=--e:\S#CH@;I_/P/NC#4Z8R+
FG^VUX_E&^B,9Q0L2SJ.A6<[D>_@(BKKV@@L4QA>Z\gH9T;^>f#[@3068I:#5J_9
0=:ZVdZZ+<JW/\WT9H>UZVb(N[T4[]0IO(f\;0J#1Z[@4L>:(0GTK=PEPW(E6FUD
ATURQJfC;/)N;?cY>A,]0cQU:D,#11FZWO^-a1c2[0T;>=N?.-K6]8&9=TVDXP0(
EGDH>Ed53c(?0]=AUUW0d-=aRU>W&OT5CEd3ZWPPR#1F77-SS[.f\US)ADfZ&dP(
?Q]D0N7SQ/3@gFd,A\.^T<,L@VZ.P80Da2+__ZPb2eA@[dbV7Y(4)6Eb]/+2?Kb<
_D:4b#VGFS-6GXUOc+7ca3S[2N(G&DTb+70/#:1>Vb^(WY^OV2:0IQ#8?)5BBW3O
^SCU45)549R&<>7GG7;2H2.(fgfab=.LW:#K,R[&.5W]>S1\)VGJ]GY4ee5&CK=@
ZQ&W=3).c,YM,W[GZ9O9d]J.6LRcc\=EL-Z3c3]1J81./1LRg]8K=KMHU1#1dIa)
Tb7&@LL2R/_8A^bU1Q6;0fQUN55Le(&=g=Ac_?B;;K4.MN6@&TH0GWTLL#<HO7;2
T,BH)H)?C3gH&3C_(VY<B?O)@[dQ+:#[b(8UeGO_a;T(&6dIYKLC@</^g,dJHM,E
.HF1ZXL@2CB<EP,R/c=HJ6)8.9FL@WU6G2P?_)4[,E-8^9d?,J(1R:bL=LfQ)DO9
4-/bV]<>EFHbKJ<P=)=Hc(>bQ[??Y6<L,I?Da[Y9#2\(LE5.ZC>FKC&KS^^@VbXZ
5^39=gBRFf)U2&(f8R1;-.Ia]LS>67[YQ:TA=>YB7LN4O8D5\I[#8F,VA[T)FES]
>(JE5TCgT;TU8/-F]=J#Y@<UT-\d474I)@<SCebUUgVg#P/S+fYTIHWA;?+c/6<3
::ZJPUKa_(H/FYP/dJK\8[APc3.QUUMZK.L6ML\]V]AL=>S(g2JW?_WCTG;.E.a0
S_8&71I;:9/Xa<[G]D8;P(SJ,eSH\H#6WIGSNc]H=V//8L_P)QI3[ANP5\2&DB3\
6Lb,&G^667_5Ya,PLV=VE,OYQb_^&b&4]2FHe6Q(cKfM)(P-YaMd]L14^)c#VDMg
0d_?G73B,G)_6Ic4J49Hg-[:=[4bcL&CU12PGO@P]:[+K:O)bZd>H02RKGGE+#78
S=?V:C-7Z(C?VL,7L_#b?38E/gO.UE]K-F[Y<2UOWQb?\ZZa+UVaPM)#@dF2C]b3
WU0]#)\gPFEd1^@F&-\KT?e;\E;\WeY(Q\EGUAP+,IZ1;?6QUG0bg9H]D_fUGafd
<.]#T#[3d.5c4:\aZ3RUe;8&26+T;8/C\Ygce>8-6;=[=-eCfM\A3<87HTeP+bL-
B<b2=[e[_[cS(==c&.)ZKO)\Z\[8&<TLL7+XS[+CE?Uf1Ua]fK8EXLL8R9+(\(@4
K-B2-3?-M[GDL(:#-A[V,?gaO35,X(55^b58\gP\\46Ta=[0GDe/S\::]H;Z2F-6
5?cbP8\Z)^?63CKYDNO:YEcLeRV\O(U)MSdKf>/P=DSC=T_afM\RG]Q>_E^G_Qbc
UDeZO:I8?_3C834]Z4#[gBXO_=f)4g@.TCfLHF3\=PZQaNH,e0gG:-dW?5F8If1C
EQ4Xd9^f\9g+FeNId0\bX6Q:(;.?.-9UW]2:EQ>bMdfP=[ggZ=8.YM6f>,A\/(H,
KaR9X1)[NaUX6VM)/AX(SMYf]65VOEUE5^(Y,[ZL<_-Uf:<T1KODKZJ-R>g1I5Z.
#NaAFA>AU]aBHf)MPJ+(IN&&M&VBec[aD0^4;eWKg8@4FIc61<HdWaRNUG]A?cN3
F8_]/9&[&4X<C]\,PGP0F<_W/Z95WHM:EUge7KI]&ddS@e8:bW0B5U(0P[LA[1,^
a<(68__CQY_&A?cZ(]J4FD^<L>KZDT6,7cNR3=)HBRf-DRe2+S>MZ;M)Q&&MEW-f
XAP5EQZTRJ@ICgb12-U@//F>3^>NYgM)\X5R4OW?GH#.-FRIKL4c9Ca1=-C/PC#d
]1+]#cgOGG=0AgH68,UT=YB8AGIaRRdF&4eN/3[=6A46=e@W>VJE5WbR2YVdXNbA
[\#&?2c\469#Q[Z<-90HJ1.cO5Q=97NS2WaF+4?J9a5Qg.0Y@?#ZOVM^O6R8Q&A=
bK9];dY+H3bLFEf@C=-d1/cXLAf?[L1Xa90<+^SKD@TDT2,/VOQF-G08=3>1>)LQ
IcFY)6J+Sd\KI91T:Q:Jd<JXA2QN>?>1N<HGKIZA0-05+_(()B5Ae42)eVE^J;cB
7)U..B;1DVb<OEN68&=3_.bb,FVQ2K58AV?[(6f^9eG).D7dK&1>fW)M/K&7C4;9
A\H=C_9f@),518@3W9E\87S42\4VfE+ecYWc,7IM\ZO1R6UCFK:RA8Yf[1DQ?VLc
-:6W4K_W/,1(Z::ROGK.6DWCcQ1Z=^(.4GY)-<R2LZB#.=VEPQeUOI-1a\27\f=Q
3CWPO[K8UOA8)MJA,SI3eNgW77eZ82+/IfB\&CS3RBaTBO2MN=T&9YUOAaF\[Q<J
2b6HJ9f3Q_,U^fK0\)8\\^&LAI@WJM\1:80;<-EF/,Td3&N5E&cY&/Ma;SO?G[QT
g9\aZ.W6SfadMI>[4\^DK,WK.@\7,X+bRb@_-SR[EA;0\]Q]->6bfC<_eP2\XgL+
--=^?FdQR:WN.GV2PU<b]fLSeF7-B]INF+ES\3&Ug)9@6(AI.B/&YV+-WZJ1/S)H
Sa@LAAgc=V9UTO#OT)U>:T0AWH(:70gBa;#Be7CO0>P)f:PSXRK[)9.MB4CV]J-=
LU0&cOM.Q8)M-TV9A+/MCDVa?TfI<&GN]X.+egO5Ud.^Mb4Je-1e@R?[4^-=&La)
Zg#I39R@\YIC=A)C&b4+5d7Y(Q?\2&Fa/2FZ7?^ebURCXD(ZcSWCZ6T8M^\H^77,
?NV#43c03)T:KN6]G&.>Z:QD,-<@>FEd/JE9.6G263K=E2,OQ#@\aO.@aPKJ#3/4
.d#1F#?Y<IZfd49fF&g<V3OYRIJ)fNJMZLB<G@80&=?#AA\#U-,##-T>RfdE0Q/_
6<[Of#<^KYFKRX7>e^S<,W3\0I64:dC@cT6R)bO+Ia?cY5143VSE)?[>,_0<]]2Y
&_\R1-:JFVYGY=);ZB/19V\CMCLAfI7Sba8A+[6G0bINgV])]1=:]RSgM(6L1W?W
+PbSV@Va0I_]UTf;PKMKb]e6C3V0B&ZV#_+.)?>+LNV.I#NWBaV4W:O0C.YGNb#d
5TfHb/&.+e],]Rg>71]F@bENX?94IGI>2[(8e,SKC#2g6:[I:6(B/c2S(E\)A&M+
cdM(Ze5:O/RYcD]NYRKaBMeE[cK:GHL=?L14W2-)dc^?M6FEFJMf@g--I@-Pd^KK
=,ed:SWf]_+d;AW9LIfHL,;ZdcSHOS5MH)/=9A6^1(Ad]39c,+XK+RE;/A2:((P]
)>)GHed7)/_>5#JY@BE5@9Kb4?d1G;2@:TgX>)A3JA6,DS:YJ(8OWA4)0T6<Z5Q5
UI)(KEDT#S,+?]Od>aMP8,[g[-Hfc?;bG]UE\QCfY-CVWIXYIT:0JA)+g_#X2Z.=
WGH..PC@5J(D8R5dRKIR)CGaDPO&2cdA?JTN#-,X/ceAKcd=(DeCYD-[5>/GH5-^
Ta[6_[Y4La/e9=RO2B4A6]2R7UN].X+]FB7.I6\[dR+(#[<:3[960>cF/[CH4D[9
>TEZJK+;&eg#SFPYSS:gdO2A=7TDJ,F2I9M+D]&4SBgCO&#XM/>Q8)VTOLY/1P88
==1LVFa[ON4I1V+,Bd+ACJ8)J\;64\LM3Y.cO(CR^99<5JBgHHUeTR<T#3VOSeXa
3X&<B-Q\^AffT/^9bJFY(->Q.\#f5+,84M#O?G_B>./b45M5UXdCbLEQSdaM7#V;
A((5F/BRJ:ZXH,<Q7U[J=e^6DAfTRN\0R0?I^,M(NY4-6L0]3BPd,?>KDKb[_)fY
0eO&AD9KRG=dP,??UNE?NU0/aC4Q.@1-fGb\]]KX6BN#S@_-BJQO9g/&A]J<&3-(
2KP#\dF_J^H^FRK1@LWfeF6YQK8>&RRLH33-\Y(T@N?IN5RXY1(D>-DQM4;>^.MU
I)Y8g@_beM-T3.#\OQMR3CNNC;A@eR..a14O>I2T]?C7_a-PS7G<]0SO/J?aRE>T
J\2C;[P>MPA;X(<fc67);?-JBC@N<)TF\QdGP9?S=TDa#8,6]KA@NcF;B-F-=@AR
O_9F4@bL6Q)c2=9K_+1Q-(7g233BHQcM[R-/MW_Y^/EG+d+,/(WN#Y2XDI7TA=PU
8;>9+F[V6/=Je=dP#A(C<=ZSLbgd@,C\HSLdC+1]\58GdF(\aQSO3cSPLI.HD,:W
NGcED\/J^ed&]7+-QRGE1#P(BNc=9TSXfD1CX18OALQ9^(FKW+M0BdC48Y>S8=A&
VF]<ACUW(d@0LCDU:BLb/4_25a[AJNA26dD^;4QL5_E#XPF_W<-FPO).2<#&4^V]
I=4D33,^<UDO=:Y.KYa[]#G(Tc1+g7eB;a-K0@X7ZcUTWU7M2?]G7>^_-N\F4))E
cE&?G8D0^.bE3#,RN/0@8K\8QgcPLcHX,^IJR+)>=V88NRQ4,)2&8T72](9AKTOe
5/dCUPM.^BbAH=eZ\7T?]RRa]_-QAcXg\P61NU+TN7,L47\IXcVH8cJ@^:K0G_>L
E:>62[,bN+DOB0N23g4?E#=CDPLYK&G4^aKW<K90eaFLOFHD#<Q07EB-QBg#,@5@
)@I=0OV3b&&5^dO5ZAa7c?Udbd7[QTTVb9@ce9@9^E\^,B3(+8L1A9YL?\4K9609
/#Z3ZaJ9^cB^738f-W3K]BS15\f>P-SfPX_/g2X(DA[Y:/A;;S54N[?=26LeQU=7
33\2)gPBE[0<P,:Y^)>MW-.1::g<06:F,HOeO_/C?G[_=T(#&cM485(0PNA6YM?C
TQ4&/#D_=DJGOgc\:(+JQU;X&=1Q.)3K9Q[e7FA\<2]0,cAe):>NF&gJU2fWD]P6
\4+T#e9P-fF>3YdJ;4]E:fP>CAXJZN5J_O#B_N]320]JFYFE#/W2IdW7M.PeF@^9
=O1Q:ZPg7BWee+6CZ+OcVV2RaI\7X06W@AfZ(#6Q[8YOVc,9bJ3#2#.Re7&=ecOW
NBJ47M8TXaJI;&;VVeZQb11G,UYAdG+8Q.GO];6BNK@)S4Ra9V/6P@g.7^W\L\87
7Ie5L;fB?;I,>O9B-.71NG&PR\L0\UfR(9aG7Ie0;>>d[bWb[_23aG;).3Vg92>?
LeL[ZV6)MTP4;+VP<-V\\2KL/LVW72PRa6_@@YR4950gKg./)UE,Kb(b#=d#dJMC
#:;IHQAI/&<^]a[RK,fJ1cQ>;7Z3-LT7>_gMc5VEWWR3b13RY9X\9;cb-19AeH\M
4fBI-Wc/1bP(Z+FH^J_)G2.H[aCSV_@fY(),<Vd>0/BDJ]O13g)baU8SPJI6:+AY
/UMGKHdT]#e/d(QTM&XZ4_2_,QBT/SR=Z6^7O_4@E9Cd?I(ZW^&eE.)=Cf&UU+1)
M\H?U65;D[?I_(J97F]DWZJ.4S0Y/.a47_:,DBJeC@a5;7O0QbUZA5A00Q>K/>]N
:7K0WQ.J+AUJK=FC^-977PWWHa9[GAH.P/_]Md+V,gPRWA_HRdF(.ZD&S)05REW&
H9]g>K1LFbc.[;c,_M?Pf=_HX00WV5=Z:+Ea+\3D27Xe1L:T)=39#G;MgV;P:IP+
OY3ZV?^V)T?U[A[X/[D&>G<F#&(#7N,#bW5G>2[ES73VZ7I,(JR=0EfU@#KC5D1=
)PVPSVc.>bQacZTREGLTZ)UGEL(MEY.H65dMTY.VC\HOF+g-9QJL5K<7)05TBfU/
?L2Z0>JOEL4[&/G0/;:P/bF\YAD6-TMI0I_J.T=YBf<cI#dA)67@Nc@BHJaCed.U
-b+c)1]KE:DI#aFeG4\=Sa,]bFV0-VQcBV8TS<QgB/]<0N=X\/Z?<1Kg3:Y;Yd^#
RT7f&=K<-gH&M?O4)OfAA<bdFM<>/CQK?2AUMXDc(&cJ5Z#ESK1;>.64@4cG)Q=Q
GZOBJg#]]MaJ(W?HbNf]YZ\gg4RQ[Z2E2SDMAY=W,3:^&_&b&O7C5dK+^8B](EA5
;@#SQZ3/.M+HE2;^ae@3QDE1]>d]?-ObT2QKX>)RI5_MBd.PAH1PfRb3=K]JP>bK
Id2]ASdG<?D>C,Yg&_3Id<XCE,e(e+a67CBTA(:7=+YQ;cSLOA^/cP>COQEFK2gc
HG>bc;VNY.F:GNg<YBL+9#@.I04H&;?Z89e_O6F[@3#e9GX#IU.gSe(+0#9K3R85
O/F>b6K=X6X&Z@L+e^#X_Q(3d2E48=Pc5(XER-V#\.;1^SbT-V7Q[&VC=>ZB&:PQ
3dN&([[.KYSZO)dADL<R_bQX4RJ/g5J8ff;(^T,5;&,+M>)fI5R(3[OHJH,>gD\d
?+<>GSPLN:D[-Yb<E1/,8U+O/&:,b9O4]1N)WVN\AQ2A3ZOD0_B?b0RT?0>X82>4
RX.<aE=Z<54H[;=M3;D(B:U+L>2,fJd-cAX+Z?T9P+UIcKJ16C=0.7;>WfQ,4JKF
a0GW2N1Ve7#^MV9WCI;@.Jb<X8YV<29..fTC54+[fM;0ZcW^XNb6SABA.PP5gAT0
.BYWSR=K4FHZ_Y>BZZ_W^=:9EC8B_&=a+I#QVYF6#g&E\R=Z#bgM^F.?Q<eP.T5D
.FW\\WJbWBR?GcN/NXRHCe5_bY0dQE>1bdCQ84+\:6RI@-/]FfTeX>WJW;XTP:M=
.]E5FOOWc0P,2?2SQ_G-_Xg3VCB=559R1+83E5_BF\Ge\KYF9HeL[W6-8?KE(B(H
]C[W#c;>gc;BS]EASM_Mb8KD&+0[g7)QGQd/QOI+I[5+1@Q>(ZI1W8];COD>c3V2
]:Y[O7?b=dB-98NNYG8/g;>S3>2U6K8E5<2CQf-a<Y>DGR:g;XHK>eX]f/C:_KcP
fFJ;f=ADQHJK^N0AC5&GL]Y#0<58bUVPCU6S4fM0fDG=U;N18?=DU0RA]f4D.R2:
D52Y/M@0Zb50[CM6@Ma&(:<^dDA7?8>EH\?ag9_94f\#(L/GJ4(OZ<_Z4N9#(BP#
MQ//[RPa+,.JT80c2c5Z>SFZ)Aa?4PNeaT\^(O]=e&/;9>)dc4CY1V;G;a&SefSb
HIWCO67QgJLX:&V\Od^^_#B?_)JU/]8=BN#O9?,cNOcBEI>TJ?SVB67UB8,(PQ9^
VeT?L/N[?fb47P7G##[Je[(V\EI1UB&gK6NR5eEV1AfUU.;GU0:F:?0USZ:0g5]C
3,V@78Q>6Ua)<N=K/X\6/[LWCYa+b8(L6EU<g=Y@CFD,gEB-(8QMF_1aG7VEU4c^
DL[WJ(ML[S?1N/:b<aU?3JM&/g7.)CRgc:6fSRGS+05bc657Y8^+a./R8aBTI/c2
I=<YG]=7N9#(T3gZ,U9ULX_3N]VTN;D92c:_XgLd::.AX?M_SUFd/g124H,ebd:^
cB#/+Q2.gPBR+\:#(MbYI8E;7cJN;@(7O?Q+.5d7:A[-b6T\>@6R_cMK>0eVST=7
>P3);K?,<HT8<T^[9..;3[B&8=4#aQWX?CI1@^aH8(VH060\dOO.cgHA4J3U<\Y]
.S?eVZRA?^N?<\96<E-/40?T]];<1FR,,6H_U::6ST[\XDFRa4a(bV@1\+C,8g@/
8:VZMA.0>(1d11@Ca4S_@&1^GX4^>I?M;HBA,E5:+_S>J_f1,5.De<[+AO:5MM5=
_A\<TL^P?J1Y#EE9)#VL5#Kc0V200747eII7Q\_+RN.O5GcK3:=Od6BJWD?M(UV3
W;,>H,cPcM.NC6d;1NI-EG((C;f0e\;LYacg6V1@8K?1/JCH13>JgFZQHEQRL-_c
MP<BZ(1QAGIeQff41T;>5HA-@\a[J:0)L&Yg0.9DVC7AAG5.[Y37Z,G/gYZ^-ETA
aKb>DZ^L3(XDK:G+:T0bW+MEK+eRR7OB8-M)R&KBG2#9d@Z8[QG(UZ8@_>A;>3)(
?,2VZFg+N9(CWT((.H+7N]Nbg?LO&(ZL.@CH<<MO7_/dFQRS_U1O;Q41&5RVD65S
9Dc^D[U(2FV1GAUQJ?<0M0C/E\-^PE-N+:1,3/0\DPAF1bGUeJ+O56R@C.A4Ja2M
/<[7I-;2</VW^0#SW)2TAPQad3,c1K)C77)?cA4XVL#[^B<QF1&cF\bVXVA+5L/<
&fYQ,5<\72dX;F&HXT3V>ZZ2YTDc71T_Je,.<#-Y,ZOO]a+M2T/-TFP3aS1X@KY^
d3?ECWfaGNLN)0Q&-X89G(9dW=YRAF]MOHY/G^O[8R+eS5X3HW&JWMGJ(H1>17c&
:MVE3RRSCV6&)4:P\g<T+gef@(>=6dW8^^:^(^.cCKaZRPa;V&/5Y[,)C]U_SE;T
f9^)PfH8KA(2AXH^<.M)=OZ9c1cZVU)EM@A8e4>NJ.8ZQa9K6#bMMGa8\_fGg>0J
X>6c?0:#<8:/OER6e=.G2<aJ#Y?(c7R\O;@1==4/Vg4eSMd&#(G9E>T)YR+PN-e+
2Y9<,>PaK_9[[[FH2>UK\W8VdT(U4g^#BTJHJ6)DHY9##9DXaV[=f^3\)N)<_2)L
,U5M;QWC][&YJP85#>3CV^S@UMO2^J>YZ]548Y,5(8-J[QJ#,G2C<@QQ#-]4-G+D
2W=6HU2R/(>+G.GIP3\T2gR]+Q[B+4C79=^(MY;KcX8bb8O9#fJE\NJXWK]aB,>-
8+2Gc:W6P2JZ7[/,+gGXSXSH^c#4g(,#ZWHcS-,(&MH,R=U3_1DTVEYT9#_6/UES
=Z^-UGNI#+^MRbO4OfN92\9bW#65HYT]?[#E,IgKQR.<2_H0\UZf(6\>&4V.^+A/
_:B93>YAKML>#ON2.HMa@Q7B\\;9J[G5WB^A+F.ecWJB[MG3D)GHf2@3c;_578C@
9QUVLK7EA\ZWd^38MUJ,;3/OJOEZQOH>UAUS#(6=OPA.9QKe9OX),JD4)C>CG2<e
6c9efa)b<WMIEIY;[TMTL>P;QLb?F4IJ;;H>JY5#@?[F2W?9)T:OAU5U4Z+K\(bW
MMZ.YAYOC/[#Y@S4G3UR=@IS]c+15?g6&)<HKXgTD;B-_0cdGR[g^?1SUYdQ4E1B
LFL??aBfE@f6FM@?&@0M9V,VECf=DZ;f@?WL+>#_B(CU^-7[G/eeTdb^C28Z[@&R
_DVU30&X5>MX2\ZUg^d1^MLB;I#V.,T&^P>=&=_B8;=\8K]dT#1E@c1FZXUeW2U2
.B)RK;/86F8T^<<1Y+DFI?NCPV^8a1R2R5<+(R#4K;N9g\1#YAgT8K:QQbC=\7g:
I__.K-G2354bTb_U]?X+7Wf-V,NAA,_IY=C#2_4K&:0g@R)<bAZ+?=QgB=>AXTT<
IBcZLDU[I7_/6FSDb-HLHJcAaZN]+V#a,K=5/R(HUc@>V3/R\@W_1I8Af?<^Dg#V
I8[C#YC=??:L/DZc(KENaB)6Bc^LWTe//.UPNO_\>,g3T4;X@_)I6e4JAY0X/6_X
2Y/5F[(/FAcLLR7,-Q;2D1VO@]Q3&^6/U>(P2(Y?6,Uc#2+@C,=Z)KQ765g&/9C6
52+E;U;,=TG5^aS=,]>VG/&P#CNEXRQ=<E+U:^&1>QUV13Ye__9,NX&fP>OV&g,(
^BU9cdDC;]Se6DGMT2FC0LNbV.<J(M3E,4Nc;Eg8]D7N(3RVY=7YW_>AA9IGVe)5
F8?U4VfDgM/U^.(Fb+gc8-1KMZ<.5aA52DSH9fedJa4g^9YTE&bW-RM,\fDb79:&
.I7C-(S.c<eG3[)Pe[K/39=M#W-CF[,0;OS+7JT5g3R3&f?#f)2&eaY>DW4gS/Td
<-J4JT-CZ83G=BPg.VKGCEbTPUc==BS7(ITc]8+I&/R]gTUTCMEEd6VTR:34,?Xc
0aDPD^0U,)H0A2YI#eJ>FR[QIfM,O_2^>01D0UM#R3]E[2.XbN0VDf+d7QSPQ4)/
69CgR\=C0LR86?\=([2g_97X&g-3PQ;P2X)S=<F98L9CGR^=@e,#\/4f\dY:-3Q)
:JY==PPM>KC_17Zf[cXW11/3)71b&EC@_CT.9AE@PE(OY\7>&,@#Z_HG0-]g2X8>
[+JHG>[+8]=W)@O(RHSGH(O\SaAQT5C^X;-f5D)c&(,T5/Q+ZHf@7>baO?O@9_5R
EV\</<?^WDBS=?)E@P_YH)J(,P1\e8/cZPE4U_R:cZ;P&,d#2fa0YLWW-R\;b+^=
F94/?eWM>6YUT4:1:CU0XVa;QOK\J[(CSeQf1&f(_Q?:M>_10W6</^I/9N@VcOC7
)b<O+[e_^WYeKLSg5eRUECJ>P/A\)+A(<QW?cfC8,20H))^C3(,e_0YC8IIgB8FU
+P5Q<29L55^];/>I=P>5WWTL4@=7]XN>e;_39Z:]=8cYRgATb3,Vb.I2@g(T;GC@
/CCBGLb^EJ&KSK]O<F^F+&FG>8TD@#^LCL44>Ue&I9-8^bI]O@(3._I1f:bUBJ=@
&N81Y4AK@BC+9C:TKF=UCAfJ5EVV/]bcQT>5)81[S_aAXC6W]CWbgYZa8gab4B[<
EdeD_NJggB[YF=C8YN.a76:2Q=20E3aLSOdbDaVLT/.VD7B_@ABLX_2ZRg\;^g20
=+6L)KgHB2P<@7,HR2;d)8ZW&SO7AaA5N0(bGGaf/dI</=F_,g_69FW<XEHTTWeK
)&8-X8/f:+V8X4W9WMb+@c2W,_UK0^F=)#cS?X@b:/AcTDQg<>1MZ6TFT;HD4TGL
2YaJ6<WfTd;PgEbLG@FfKT;fM+;;cd79XYg.7d_f5IXbQ?&N2_5<E@(07]SX([X7
&RPgIQd1ePTcVKJ)aWGDL.).KF4H[g+-:eB5[0N#ge?]Dc#e5e)aDW)39KPW\Y2E
SUT&\.L;8.0aTdNBXOJ#MgE)GJ<_L@6G>:[&eWVCXVJc+<_4(N/7G1[58MKSO<#A
X6c/^>(1E.aBL9daI]0(/d&9?M=;6K^Yb#Uf#U]4M4XNW24HB&.7YR1Z<[Q]I=;g
)T+/0LeVgSQ(C\Aa&L:I@5/5YE:Ha/O7DNJ(3IE=7X5GDQ5^H;-fL/\WTH.4X8D+
--L0<dPPbS:WX;dG:0#G@PfW&IUIQ&WPR6&2T_)=Q=DFdL=M:95Y,?E2IB[S5?\1
;SeX/HfX?GeFTE.AISe43ML:J#3?<U1&-_E\1G&\\,cW&1IJ674#/OSE4_M.=X(F
^g?9.P^;M:H3e[1UJ:-eK51@Z3b+TS6U<5.YVI/d/,eN3UfU4K]I8^G,Q-#;U[J^
I5;Rd[IaTHc29=cXVH9D[A,cIAMBTA8RIEf5D^a7g-DP+OT(+EGS(?>N-2(b\<X#
3OD9^]E=(&5;WAV@H#1,.7\;bM)gJ:AZZ^cG#S\\;WVM4L/aU?&R=8WZ)EQ;?V7L
Y40gg#R8K@9;OcdP4Z?1Y([83DN^_E]fJ1OF8cX84(L&\LXL).:c-ULEZ\WO:6eB
CMAOZ(4b\AXLe_MDcNR\&CF3[c,+RKG:ge&+ELIN+LTLD(U[e:AI01XDOOc7)/I/
^49OG95E6a/)?7SLV1KL\44TI\12KbHbS[C+>_C6-KJM^D8:0[gcH3YgbVaH86/0
S=)c<H0cH[UWcMV;SK9(\3#36QcTA,2cABEc?GAe/4F1##/+ZQLJ&D.:-\YfPC>L
-gU,6S/OeHA6;B.J4A>JW[gcY36bf-EF>c1)_Tf:g-<eaA:V6_<R#7>MJaXE8\84
QD0J=ROQeWb4JP4\MRYBKUZA7/#M6N(8C]#ePf]Z#09LRJBP+85MZ85:F@R9K,^H
]<Tf9+\1V)@QAd:bed9AV-eFN;bOZ-U5=G-25GOH>ZaYKSU^/Ia7W;KO2T7QF;Y9
4BE>cXT+DZY8Z5ZC+LJbCBGUJd.F51ZdDWXPVIgVd+1.Y>1?3.8#DS..F322&F@O
;G33_=8g\4E7I(T(U5dd3<A7g5UKL)64eb5YgUSZ]g31P(_8gFZPfe-BTe@K?eB(
GdAR67P,<>R(?5RMR@b4Z=HZ6d4XOVbcC7:G<WDAVX3EA8L?S,cH=F]Q,,\I1/gC
Q4<8L7J[;_9B=dZ(:=CeJ7BTJ[gX[EUE=1LYP)X.\XWBeFI);\+QgOcP)D@>?>g<
OV@\A(GfE]A0:&8?.C2?PF#).[a7<RQX#9b>;9AEM8(=NFT9R@AdRZ>5O,=Lde(]
_&AOK8E/RFEN&Gc/K[644)N2^3G&<-gbb5VT/T>](-/U;NY,VMBKJPd3)_L1_S#J
,&X>1KOXE=[^4NeZ)Kd06Ug>I&WgX=@OE_DRE-PbJ]\d)?]Ra>b71X(864&\R/&Q
AOK2JfNO;1^e7CGY=>2GVCXBT1SS(XgC9C]bPUAFZ#aMbJ5FP>.CTB@LSfTdD)UY
Z2R]8L,]D]YUQ#.fF;39GF21Z;/]EUB^K#Pf:N#HfE147OBMN2\#F.-A;0VAYZL5
eWf;#BgF0Y[[0P5OgCEg:;]H0YU5HPG&#NHUF=V=]47KeBPJT7LIYWH#+UY=U+-X
Tg)bTM?GPaG@F4[gLA(1M;B,OB;S5^6Q9_(Kb9]^PN<?6Qd>3U\]?)OV+f&)OLHe
(N@/(97T9(@6NG)FbELB8Z;T5Q=-6X?IfR&g@]MU(]d]OB9&E5GTgG2&(,:F^<gX
,O75[+GP\EMYDLVF3g9G?Q</0P@NZR#f5VJ4KSD<(A?H_/Y]Na4Q+bT@<3;A+O2G
AeEL^\&\^&2eBJSbCaB1#6JRP7KVd15)B6+O.2d)g\S]Y>:EcT4Y>QP=N:^eXW:c
G2-7A(WL7.KB3+GcY0^-FFTE?LdPPeBMSWTF4+e\N#OX:4\cUb4+RH+09.><YVEd
d?Sf9NN^c,<f(cY(EFQ]5#Bf5F(-]?WG<UUBBd2gZc)7W[gG#,N77Y@J8U(C;:I6
,]^ZD-&;-B<F>#?1)WK8(_]IS6&b-@0PC)2C=3/IXY^JJV&#>]S01bLBHCT1,6)V
<)86>Hbg1O#Tf4?_FgVVYVK#Z#EL:K+P;SND==dW?=7J-JR\eG:UB=\+S>FgbC]5
85RU294K,@G-C^-TT+9I(ATFUR-<3(:a097@eEB;[H->HFM#4HSDeP&d,)#U4MT5
#M9;SLKC75NSBf\GN-fE-:aCSTNS>V_G]EdA=Y6eZ(KJ9;U^N=XdId;HZ&7L#(S\
T&QQ)O\7e:6U,,9Pg;eJJ#OfFL43E,,8YWOC^8JRMCId8(4/]FBP+/9fQbO:<BM-
b[;gR#6&81gg7EL^1U(Y]Qb[DHG09,g5E,_b->7\[a5)6g(J^^0IBO_-S6d9ScPe
<EU6&T;;G9L<(dfbRdY]0]7.J&BMgEBEKgTFZ2,fQHYDcIb7\B,HU1W.DZBf<3JL
AK>^g&Xe2GF1cZ],<^PdBO?KM]E/ZR[<8QG]#A1XJ1bg(W],O&,R9QVR@4KZT3J[
:?#De5;WSRMS-W04_(\If-R=c_+\E^R3\_L12ED-DCQQ:=)&9J7e>0CJ&bA15:(\
dD&YN7Qd7-g\PeU?U9G:[YS(X4N(b-E\^/Z]\^DFM-?WXaX2LdYM-RPZcV4R-1@e
#NbVK)Z(+HKC)JAC?84gHE@<S5BafH@N,]&a@I3;JT0+C(/E,Y]>[Y@^.NQg]fE9
&XV6\H2KGE_AKbTNM_:FH\9f(;ORA>MXKM-?1PM(6Q2\G&Q)g:,.WY4-]Z/C]KBV
IG#S)X-T_6?GG&CQL26>8UeeP+R8EF(1F\Z)^+SeK_,&c=F^ObCP[40H[A.M6YHK
d]O35f(ZB[f>WRVaVDW^JgSFU;H<e[e]78)c<HQ-7/bRGOf>>HS75=@.2>UeUbKT
AB8EJ6?@+abNfJ(^+dQVaYZ>/=Z1\>PG=]SL/.+RV<H->BDX3#SHUfB/-^;(01=Y
X;D&&T[KEHSA_Z1a)c^>T:HC)R@TA,38N05;M46@@SX0UL<Qf#5RV)C,D>JT2ID-
WO[FRE?bb[VC^D?g1GZ#ebRVMFW(V?.@DF[-A6ACAT7+[A3OY_\R@H1G<]U0Ge3I
5[Z3H7BJ(2e<?V4K57WFBe1Ra[DAQNTNd=Z?/S.a0<D[&D^,]daN6e<\/NZ45OEH
?]6#6C+,&))/X7,a64MO#_G>bK&@;#PNDKRE[LHCA)0>Qbc6R9#fKR8\ADg5DUY<
;XQLW_:=L#V(A655_Z:Z#TdEX+>?d:2)U_[U:b):GV&\)Ma7Hb5P78O292VH<1]e
HA4Z/3T+_8J]WL52JaIKNS8<./3e=J,3X/,20LK;6dZ9FCc@)bg2cU>9H-HPN@WX
fJc-L,PeQ8G/#4dI-1KV[e,91bYMG<AWJSg6&@^V?Q+8\ebYYZ;3>HT/HU5&,aSZ
;D4@04.Y^W\?1;;&<2)KG@IBgf;B+FB2/2_Xb;<,35>CJ(4f<L-2aSg8Z(6V)0WD
J5SB0(FZU6cK0+De:aYVYJ;7fBFNK^[L[[9c_W3@3L066X8Z7?C(][)#L@e_J)M5
5MI8W^O3Q,L^QFdQKA+b?L06MT8eHF#EdP:23&.cA#?8?a>R:d.RfWHA0-#55dH&
U5&>)OR7JTW&I82=-bR?IWN)L&+4>D4Q2&fV6JS5WY-S)L1)/MA9:?I#N&Hb(:+Z
OP29&f#((<\4Z:AgF7EHVGf6L,-PRPJ5QWGEbX/)RIQ;:..8KKNN)K1NN+g2L/BE
9.?YfM>A,XPQL6ZFAMUYd>gZ)KC4YcQ#+/-4G_4=LOA>__PBY5N-e]74RM+2QAJZ
GAXZ3YeY06OecI0AKPcH>J7dM@8a8_0WM9R.MIPY)4Zec7Jda,:3B?Ead/LY)9d_
=#TdP@0NBC+-=5#U5C/]T^]1JDL2MDI.g8<f_\H++P6@#NX3.#Z<^2fbHACg#b@>
XMbXBG;PFdZ/dfN&^]FJ4b<)UZ75M/3S.=.]=-Q<=QQI;9Y,2d+TJX[aFTC5G9T1
2LYS/-LH1Q=Bg#J6&ZM?=J5g^@#DdddU_XH.2ZJ/Bf4C7TM[T\U6P/U9I,\-Y+g<
##S6:aHd.6#;K<GOWf?A/E/5bG,9^]T(P5<CeD>FAc3Z4V4HAU7gFg0XgF<4[OfG
,53;Y28M8G.;:?&d_V0U[RBEK@G8?(Mg:QB9:_;+X02Y[^<[\QGR3>9CAcKb)DGT
9[BVdf5Me7eD@e6X<I03D=NNB;55/IX1OK\@>,S9J#L7SP8a\f18R4OJ00=B@eC2
_Y<Af].\D/6dBdKL>#-:JW^V:_+[@,dN@-.6;8F-d:W,IW&3EF0Ze)(VK7bf[g]9
O9#Ze><Me>(U<<[HedV?]0YB>[SMHPLa&Q;b(P3OaZEHMaLdQ?f#GCe8JfaAPLcI
QaXgP)1b/G5V=FJ]S7?)JRPb&D&=8Vc6EffOWFgZJ.NI]c.6-G,.D?,),d1][N(d
ECe8g:Y4B8\^(EH:\g,.bT@gB=LW-G5Y-JC[5b7F6dXRADY\/)UE^HC+fYV+UJZe
EPUAB9DgT1SYgYLf1@H5A^7[XZ2Z13d^FZ@.@+gTSK5A\TTQ^_3W84+.H5@T,[Bd
Y4UYL5IH.bg=.4/)B4P_<>Q2fe2C<LCWY;E56+CFHX)=D;aMDZ=@S&ZBT0QVG\H+
a9KU?<Q.ARR.AD(/W9JDE5aR77/7bHWe1-R]C?a]2)48YS1:[0/UM.b=Z\YY&BV)
@/X5J98TIGX:E;:<Kg@N(C4B9eJZ8cGd5]I&0AJEFNEb1?@c#(+XC0L8?21GdMCW
4]3dJL3#2b_@,0>ebd.?f1>2#?5UJX5VN0I&g<38E9faM3>5BSE@UA/&5JGKJP(8
SPBM)bUD7V1d(f.S9&T(@L]0b1>,<W)[5E2&_=ZDN9Q7#G+Z[BbX/N1SO/B;e<#D
L5#.:-EOGAAD)5[37f&]4;dZ96;01<ZQgJ/SZH[>d[D;TTHL4J)fL4a/BcHY.G^9
MYPUFXJP:;(1;7+1F0bJ[d6BcaR-B(7MQ][RWa;H9gEA/d7STZ6aD/ZX?&Wc=\[X
K6)\T(Y6d&]QJIDLHGK6:HFMCA7C&4JfV]#fC-,N.WIf549W?]73+E^b,e>UK;E7
UdG>/[;be+]2]NRRB::=fQ53fA4TWEGQLf&L:AF=+agMTTLTde.-S]I>V5JU:P?+
f5R2^(H+?LPI8gb7Ha1WS<c&HKBBCa/c88,eUO)K<<S[=Md_R5.Gd+)+/VCKffDE
\X=^&bZb_\FEEY=3UI0aI&PX-6G^LB4eC#T&9B<T@N-a4?1DIea62+f=GT-0?H3-
L8.(;\SUcS]N>&2]0-,T9=6ZY0A_:EXEAJWQ,9YM9034>APfKP1bWW_NLTdV?IbF
8KVET@JAE<NH25:,<:;90MR3(FXV\V0B.F,C[bSCbM+@<R7U_0/O]EV0O&@Ug+JL
^R^EI+T=LT44PW<#92-<C+)+]A^Kc:>.:J;A;ZYZ@5,L#MK)Q^&.5+)RO<SM2F+>
O-;<:HdU8???26.43;-V3=S79@-f3A1cBb-dgR/-)H:(SdVNB&JdBG>b+Tg;]MM=
GJJ<IL0=d)#):_e7<.=WG-V#NQQ]PK]XA#I@GUS#Aa2GT<]1a;Q5]Le]/79[H(09
2&+,MJON6e,<MB92&-M^ScEf6+7_C8ABE:cSeI>ID02=LT./15L-@Bd=RX^(.?gD
G]_Vd2Q/Y.VVU:&E]+aJcL^A5=T-E9(K\TUG0U+V^Kd=(>#29C@+cZc-cFE:(-5#
3@9C#BR>K\a+5W;>b&K6N3e@0E]aAMJB9JXLg/Q2C7=g:0E>bQ#@^1&<gKCG771#
>I8H?99V:gdg3^_Y@a[BFNQDbZAdQLdg-\4>9N_Ed/d==BJ4A=aPdHf=@VdJVP(.
5J:QIgX)G&T8L.aGV#)QNe0/Nc1g_]J6UV[ZI8.gQaK[JRO4AU>4_L5+H8-2=LcF
g@7&I2\(fI.9F^NI?.&#5),0>+TZd9Q:Z-RQY.=3E6<Cf/,d:gXP4e3,O.^b^>]+
GDVg0U^@DK=,fHCIM?[340<^caEL.RWeeaeO7d1ac7(15&Z09Y7&4:2,L#<VNcOO
;+.)-V:A-(@g0Ue3T\;W?L+TDE^R5e=E/>KgHLUCQS<=;T;H)GY+)-\T9RCS/.[A
8S<MT?QKE,\)#5Y^1I4\Yd9(+-3R.WeYfN,X:N9=9/NSF^gTWV30KMa68bgYUED=
@>LJ81;I#H&K(fE-X2/;F?KGAD\H,+3M4#bg((3L(XY^7KD#T(_g:^718N]8KX8B
2Y(-(g69-BA_A>He7DM6#8G#b>M\O(XLb8R]ZV880G?S9OE9>FJ4I9Y5@:g8PEd8
EZ&2MeQfT0fO,ASFMG,=7Ub^JYe.>HOVG=f@dfc6[YHNfcKg@/.:U-^L,_TV//;X
_>]4K@M@:>)9L&-ABC7-W)gM@ROE^CYeO]ZI5C&I4UQ8:G&HB2-W_JCB00XITI:g
.+,UWQb4&a:@Q6EAHBb^+(?I<ZdcVNGKV?,6;<0YdI^@O<B0M;\X)^=7E[K2.7S.
60F,<@NL2++B:#aBIa2IVP[R<Y#:.ST6Cg+3(8#d6>BWe>6;48PHGA;1ZC^SB(I\
M3R__BZX4g>59281RYH@,Bg4B0@N>P#_N(DGMR53?c#BdP4O+2MF4O+[Qe>\VH>e
c^Mg]/f1B5/bb1cAdQRPL#Z8g4W7)P5SB9W,f0]A;NDNHG-3ZbS6cQ3+W-Y#[S9F
D+eG1)9;Y?/JE#FCgN.<Y#+(LOO-+3/I1=]a+aWL+LE1]eG3U&1_HeMX;_&)Ga&5
gbV#_X0=g?ZfPONd3#\YK&C]Q34-FW#fDJ<<->VgU00gE=fO.&]\5V+Z^R/;I4IX
84I:EaP[1)c(YL6TZ])A[gS>bWZQa/J3X)5,5cGg/DLQ)B7F6W@N65VDA-GAU:I]
[GO4JSf1CZW\?Qe9LPfdH,g>LC<[\QR,a3H;^-gCA<0UA5[+X]2J=H36;8H&3)[3
V2[_?>TLbENf<5UH]4[/eBSe4I<Ee,MO-e22>Nf?Fg65Z8@[(F<G3Z4=^8Y6#-M?
]JN7cOP^fDVd>gfXM2G5?2T#S=[a_^IW\&36=H@?D>Uf4(GT.YJRZ9Kg,?K=UT0M
(Gb1dLa4.:+<@RC:(0cQS:d_^@g\?I[;<Z_.OT/R8:/69,&([ESBK,[J,UPN^M+S
)QYVPP2NCGKI3fXP6TTNQeHgHa@C#TH)ObXfS^?K+UU(=6HCWS3F)6BP/X_@)9/a
,Q;L=4]O8CKSfU7Q-+OJ3Ce,&40C>OPWWR(g\L;TR/,ecQgN#ZZ20AJP9M/Hb_Pa
(:G5Y,7/#8B/^eIA:dB8A=QN0P=1((T^d;bZD,QT[M[E-LM?1_3_QE&BEe4-I\3N
=.SA0-HG=BZg,6LaO;IF[f^^]>)A_W7)dX_Y#b,,@\O^Y]:OAM-TfH:5;MH@AcVW
MUDK<CL(D:0T[W<;>:]&SCLIAW@,DXL#T:Y\;\(=F1V.d#RM&CVeSQYTD41VMXSQ
.-WR54KbY,3faQSf4A89Sd&VUH^M0SK.3\JE/a/<)D/>J+\WG:+>gSAF]ZP-Uaa&
7<9&0a+V<EY&425-c>)>FVWEZJPAOg/K<<2c6,9a3M5gcVC&O@78S^fG46.,NDH8
c-8YLAH][VBMegE,6LJIIW>Cf5I/@3R,6NX],7b+0G8/(YdIKXd+[2)UC]Y<-,Z?
RRAfga?VS@faRAJd=[TX+bYD/P9<JO/7-0B[UKY&8^SMZO?LcK^-FG?8,;0YQ?IK
/4WfW]3_WKDgDY<E>(G4LBPU2b>XL)?9Y2KRQ&4ZZQP7S[/?WSbfXAB=8VcV>A3J
X#4^XEK/E2d[W_F)+5MFR#KRA/)8a39Da6H:9RIQ-:a),KJW-\d+dBE8,7;H[?HY
:P,-E]JT_+gdQac)HOHJ(+0A@I.(a1c1MGFL](NP#@e6^?)g7N[WPCL3YdD_GKDH
e^dML.)J#M#c90(NPHOD558Pc9ITTB=A1d[&&aTIS@NRP,&_fE5d#eaX0/\O?QL;
A)VTJZ03AOUN-<KUR4B@)K_H[1b4gA;5AO]12L\0-eP.NPZT<Y?VA26UNU@L@PFM
:<F;]?ZO\([cB^K++/HDeX,4_8K]<Qf:HJC]P6+F>)=KNNSA8][UD;7W>=?I/4Kg
?;94.MaVAYKfY@K81->GDF@C_,5=_&XFF]+6VW5:P3SK]9c[K9c#1]d1H)PTSaA2
g)XL5..Hc\^&8\7f&=K/d\I]^TLe+\aU;+_I04.:.I#Q64.P@&#\b<F^N=G,]ML]
EfSXB,QO.W8Ig\0,V.(N-+SU0+d)<YRN.=gZXDdcT;,#K<KB7B.RZU.gcB/.M<(B
<D:e93?-KMWf=,5d\b,3O(T)9(M),faGDV#<AV2&)QQ)&Ee6^NXG\YQV3/JL_;\Q
IB/+>b^GbR0U\GE0FP/.KZQ.^H;BBQ[:,A6_1eY+/<3.7PJ_23?K,aI)AN--)3>?
7:LN:ZV+4SPaO1\GBDYJ:OWg4U=>7SV<;^aC@FQ^P4LJC,/F=[RI7_QBY7^a3bZ5
]1RYDT(8Y4RW;c62g^)Q7G,.8FS<f04NaXQC&Jf<Z(PX6(e7,T\cc(H#DS^QB@FP
>CfgOY#0^PMFU1;U8RH9XVDKZ91NOeYV\dA5ZeFNb;7@4.Q6#MbQ16,\44<8,&[K
Lc_Q5Va[d_&C35)QC<QNC6dO+:\J3;P=@BJEX-P\8JK-G^b+=<Z::A/LHg=W2Xb,
+8EL=@G3HKNga(,(X&0@R+X_2b[VdfY;4,H(64G^:eBTU)G0/Z&BfPH4YSIT,.\S
B7afV&VO)H_98DF<NL1B=<3E.-4:7Ce7fSGJgJX7DbDF;dD.Y^+8G_==]/6eddf+
,R<VL)DbP=a4P(AY7<6:<:&/=^&P+e;?ScBO2beOfX8Ce33;>@0ETR&2OG_b4M8S
N\)a@E(=7JS)]1-]6VJSgTCMVH.@F2)QB)gKHYbN0fXHQ0LKWBP<g[2?=3,#X:R:
FK354O5M=(aC:_BS5&SOF/eD-&]b,RY)<K9Tcc1KV]1a_?2+a30^^ZVg#]FPd5,:
)L<_3U.df(B)(#eMB.Kg-_17V);:O>d/&ZbE.?<@gfaXEf2=C4URBK@QQR/_RCXR
&<OGc^2NeAfXD>FCF=WF^f(-]QRDBdd(-9@,TM?-2-RX4@CL.b;=9\#\5#X86(W@
Bd[]1^TP_3,VO7)KF?Cb-).aEec?;Z9[O7__>ABe/A-:9K?LD\c\45>0_)dJH&H3
,?^V26V45\EbYfD17]9:8)5+9d,U06QOMFJB^e:R39f_)g](d7Y2F-NTe=;4=CU&
/12BYXg>IJQHfPC_FFT0UeP?MJYeaTf)3d>7[ANYc0+a0dLWG=-Z+.L6gGVB=2[E
:MV.-SF1LC54Ig;Z664?Da@YG7@YRB)Ddf/@4S9(SNEJ\K9E[>+dK]+47Zc[8:MD
Vf4^@#9:.bX-V^;,>03RNg(#SC@:X9XZJH?33f/>Z)aZGXP]=)TS()HM:R19_@JI
]2-3V?b9;L5N6_B>OSTA_5KP>8Q;>#A;@#O7Nd?\O,)VVgK2)D-Qa7EHW:^(X^57
+]d5^J8(B?A?R7D/0RXYBc2\CEg=->+Z8=07aTCUHQEXE0G]#O;A@O4Q&_G5[-H&
aBTM0gM6eJ=GDQD1g,AF;?c2JW\L9<5]NAcUG4c4Sf_]YV)8dSa0MW\H95.XDdDb
8\DIcBg[KS-C8[PH/_/?6#[]e2T-WEH>)(eIg3]=G=(W&]#gWBbUJYB2]\4\;^32
5Q=@>KZ1-\E=F:c]^CZO:-GK6W4LRF^ZL4GSZ2C:LLV/LPJR3DL4:@9ULc;8S,/e
L_5#^B4g?_>7<.R(;WRCb#?YQe6XYaKLcZ;=5PG)Z8GVYg1b.Sg+>_dP+E(J#O#@
,@(:TTZ_,>_1B#gT2-IFfeaW0=[^T8KW=.GdJ_.03?f0EQ/\U7DQcPg_6a)/7+V1
3W&K@Yb_##1EC]R,>&#8d@_^-Q5U&#UaC8B0_F&@R,?@eE:)GSN@+?Y_Nf2/f)BQ
?_;6MAaI?KdI.]<\<)5?U+1820\U13D:4OB8;a+90MV)E9N2d1(I@M83Fgda)W?@
=c(=T[8J+T7<F2H_f;FZ?AHKVH@>(J@acB9#W&YASS[5;N?eAUa8:UbQU.FK8]/E
9<,U9BM]e&4.VCJ&a,9.+25-\fQ27@W)dcS/Z.6b20B<.H;(@,)TG[0W>+gfadYD
C?dab^[[U;8d18^MVOYR+Y2^^;W-XW4(K?XBS9AP<RJ?/6\>#AdDL?&#9NP#)ZLB
#@5EAUJd>Nb=2LP;4O5TD-B1ZZ5O34<bN7N0+PS)BQ<@=D8B+ZLKLc&V6BB2[K2S
ecK)EYPU^SF>C1#7GPPb.g7VgX@XHSXJ[95d89BC?#TLLDF?)L2F01HR,C[O(7?(
U>X)B?g\-?3ALAR]e+Cg;H,_2Y_.A48QNAf:3AcKVO#D7JUC_+)d>9UI;EA+X-LD
PXP9X:a&+;>B\HYF</Wgd3LEb+>./N\R[]KgCQMMSHS93R2PQ5[07[G9dbTO_,G<
aSL-+]BR[e<bNbB6J:L+L0+NH6O2MB89R-)]M].D7>_IgF6BGECN5KV/(Ng)<<@;
dEf@4QNGHS@TB]V_\,.]5_R<cBbYO5-<@5&cTHX4#58B3V^;J^?0P3>fgTa6TQ>6
X1.G(L=#(]:D@Q.)<b\ZN74]YG6)L/#D3^:]-0N,(U@fQ/GNcET23d45>>^<#Q.2
fT@3;SFd0W4DRW2VLZK\9XZ5OR&-E09C?]._B<Xb3E)CXA:fea7D@J0Y):KaY_CA
,<S9b#>eMFMGUG(c1a_UP6f]T9];SDO4Y=M_a8UDD,cY[\+0Z(ZH5G1P2B53C+=2
M1f/-(?R]ZVG)G8T(8DAH424H9e/BDf]?989f-]f+C12KY_f4PHO^.VdCbE:MHV+
R1HN\3eZ<(R@@_B\U\H@C3B?2(1EZ3_8+8;@?aTC]J7d]]\I.3\I5LJL[;^;Ca^J
4@-Z:])Q-]bK&.DZJ&A-8d366OEg&U2&+Jd.&T7.Na[Gdb[>Y3#,J?RN1aC&\O5-
=[4RcU[[YP8f-H<&2,&K=YCReI(bbQbOY&3PU43U[aJ=XJH>a/1-3.EXOF-@+B-f
Q=)O_f]>+HF@XG&\--X?=AZ?L7QB7L.-N+P@Z[,GI[AJb+4(5LW09aM3JYRAZ-ab
@c=W]BB1g(A>T.);Z<1MX>5He;(O]P9aE/C9^bKH8/d:E77KMM]YQB=/0#:c.J?<
;XB_<[3-R#_@:cJ/72cOSV(0\2:KHWK#.O9BQ=fGOC0O&P#d&#98-(P?E6/TN\T+
2URI&=U)5?,^O8L/]30AH,HN74\Q?-:?.9MX62]<_K;d+:=2UI?E.??]/==H90>d
L&IQ^19=@,WZ)E6<O2GgDb&@_aU[0?=b0QEa]g(OO=DV@f5L4^A&B2)A89UbL)g[
767Ee3B0XZJ+VceQ_>Xb9;&YS171a;f_+Xf[K1?EGC5/GLb/f(E01Sc8W7d8A_X=
27TC(,eG+1^X.g(ORc7]CcJ2F0:3NcW1G)V..C26Z0E4,g2K+aHH^5.Q9-L7,M0<
]d;3H?UIGLdDYSe2>KeV9L7L8)Z=bCg&1gYW3(#TZUQW3_^A\Kb/JbK(9H>&4H;e
MTFL2&Fc/QODgeaP3OB43[6Y<Y@I/L7=]C;d#b]fY._B)2(XL60T56d^?KWeEb^B
#I]&3a^,JScGG7=<AIJJ0;eB5WTBX:MFF\1_PT>Af&M@e,I.;\4E=>+QQbE<-8G_
[\J[+Q[58^[V_(#5)(X>41;EUN=fZD&Y:X0O.:W3E2:/(aXWg;UBecIDVfXS@J21
,S45M]KQ9&B+T(P79M]JUAGE&JY_;g9Cb<O3A>\L7MC3.AC/8@8XTESeKXWfLA+G
Z/FeQ?LfF:(BXS305?1@fQT36@UWS))I?44\J<#ZA<-c^Z0^=;,FHLH=5EHY6B9S
Q9CORD<&G^,YcK=<MTXL?KRIGWB7OUb]:DC2I3]bDVg4#98K9N.AeD(5:;/]Ib4A
6@-YKKF<NXfSQ,S?c,L,Y^K>E:7ARS&M9MJ@^0RH7GI@4Qafa7,#\+210;T/]cRW
Ig_RVD\_4067Z\3/K-0E5SNO&B&_)OUJ=^D0?+O_7VKNH-9\.Y#BTgMJF\Te&PO<
^11KI>&)60X,\[)#BJe)ML7G;QS1?+ZM.dZ5f#=>J1)G;Z0MAQJ@2DI+#Qba-H;4
1400&-[#eLe2Pf+@C\VaVHYd0dGNed2IUO4R?0)NaMK;JX[SAO:U9TFPaUYX(3fF
]f[=cP_JWL2Ee.^-6=SAXPWa6XUCM^9F\.--=L-SIec_I_L513)@WK\.d&&&4NQD
gUG>D52L]bKV&B:KGNOZU_&F0(J[15,GM>aB-)8<?2MPHJ(BW1LNN.#H/9[KL]4C
L,[XJ-&4RfPNMK<3F#1>=O]A)]P7XA=ZK]WTOP7Nc?C-9.ac9L-Hc2fIeF;5?A2@
Bc0PK]eA@S\)Vg1gBR1Q1Z@c/Z\D@STC/G=06R<]H^M@^>1OAc:a,.?T^_+C/LE,
@U#-#@PV)P>MZ662#Hd7,SJRSVOZ@MU9;-#8HKN+W4&O&GGKb106EL=IT@4><3HU
PE/deM:4SgW4(/#JCU1359/\8^e]D@O+.)cKE/M+T2EcFP_-+X#cE6:_/M4#Td0[
&3I8d<LS5,][)^W^dUa+^:X?4G9Y,2Q,,ENCV7K5bZA6.IJ2).>SB4/U3L9+)eT8
WMW;_M<-YZgf[aEJ<YW4c+5GN96XSV,R/@WA_)=ge=@Y+NNe-YQ]bZ#CSL1]C;UM
]W7;5g@9W5&=^C6cGY@dU<@28f<CGN9W6Df48XYQI8WfB_XG2aZVKbO(/^3aPH1<
I-Z23D3M7UGFf_PK@#C]b#<,AP>0J7a>\K1=]\9Z15gXb2J^(N70\N7a+/#:V:/,
&>#/U]JXF@D+7_(B.P^PTDP&c#[K^@c&)e)VC5[MJWC,<R-#6QZ?4I=L&DKY-2F5
&-@Ig.AAQ65>fM)R^)HT[CfVHE_.PM(PCSXXD=>D)HVFb=1+99[eJAHISB?FgaRI
:KLY8.F6;&C)56V)6bTJ)7AUYFFJ]aCb2;[DJBf8J7JL_[e/1]K[5JB[Q)R,cN6_
GFfZ_,>;g@2+,\fcg;9fEUOOUY^5L-1FCbBSBa[6(>.Hg?UGdPMLU5(g^ef#UW,=
c]EK?@:I2CX1b;#\=BI:8-Rd78K/6#1MEO^YD^][Q^90X&>f3,5/)EMBYIDa?>#+
.dSTU5A1XfKP;e&g9?+TPZ\+:+C3KK+/a0SI2b3_55I_C,O#U7T@/>f?=b\MbTT^
?D0W\GeGLFSX)0f>RGc@W4AVg#aEg.WFe^<1;7XQI>BDBJ[a\PQRRWGgLX<#.Z]3
c[??[a)47#(X5X#D:/[WT4A6_],\.9&/+.MHX-6B,RC)<Q=f4>aS=&gdBPcY^W\)
\,DX^VQN>V;I>WaU6fQ7BW\]@6&P.:^gHdJ8,Rd02ERB<+_.N@6S0dUZNb#Ig[2/
^,\LT:I3_=1AHd+0<=,X4aIebZ5K^G2/\YaVg&aX5#f.(6Y.5F^fY4b[(Td?@ZN+
c=@;Bc)\Q=fC<^0@I+##=+APXJ3:F2?g<B?e()<@@OTbQTeHSILQ9TQG]=g&F21U
0T/Ee.(?5WV[74-:[^M;T+G??JH:K0/PS:C++eQ:NcVUT;Uc^GT0RD7D@S:>>AZQ
Y)@QJ+7-6.Y,):3P^g[;5:OB^[PS/_dQ.aO6FW[b#6>5,[-_>9O@,cP]bI:F9F=>
#3Q/=ePe>+>I26LV;X>+)f;8]BTZdH79M6OdUHK?;\?P-/Y,OGV7:K2-g;5dC4f.
;e1/EQA_cN\34KJd?6;V<<^E0cLIVZ0ZdT22<=^2A#R-48H?31fF>AMQ/Y]ac4V<
0;fg3bK\4CbN5TNe39CfW/JVB&RE3R\CT..99IW..M/?U\R?5_;X-Wf(P.EK7K2[
g&QFC6JBAV2[a7R=e::L6:AJ\&Z:+N]7)1S7P?G0][\.>J8]7E1P[O4F>M0V34;/
OTYgJ_PN,RBQQVg&:Q3;94V06<?Z7+=\2\3L&N_aKV(A8YQa3gV[)IeT3e75XK55
Re6aVHV[Cgag#>&5PKEDA6[,\S):6(:MaKJ0S\3C>55-^V7#+<bPS5IL3V]GO?Q(
8;F;UZGPe6J7GWC2GXN[HV>a#]c@RVb,?eJ01=PWa3eAI>G=BI5#c\?D)[<ee:Gd
GLWZ.=U^QIb:MIW>XO/@Eg_.><O#cT&#7B3>@Ee168;fd05M^FR>VIe&@J6RVNJP
E^9@08#W\P9f##WW4fS8N#]GTKdbP<0IF<eaS1(M.<J5;BV]NER7ScKPU[KC9dF0
WTLe4C]3R\c=+ZaD)HDS[=;3JF&OG;PSK#S:F[d\;gA&3=SY&&^C?\TLOOX3Mc::
GDPF(KB?585>JINIR=F)B[U.M_PH<fGM>3)C5Icab5]EaJ<NA0_C#Q;IR=E1XEfD
WZ?5AX7^WCfZ&2b6V<9S(TS=4ICB7V\cgMcFf1;9;4<9?V52#(?(U\UIEWE^N0<Q
c]R=[GR.^edJNbA>2E7&JNegWY2^_TEKeW8GAG\-&S.4@C>aAeS]9RcIWU)U>NW:
R?//R>JMd)DWA0CED&-NO(5;GPf;2f6Ia6QF1]A@d\AEZM+FF&BCO@#OPYDDIGLC
Z-[JKQ5Df&]:8-T^6WM6G4MAeCTY)SYdA^3U2^1AIfa[.FFF/_AN4\+>2LTU\#.(
RQ:Wcf#QZJ1V<2HJ6<,];+5=-e[8NK[;C&8QA:cQC8<Z_V=0],O,(F_V?MaFW3?D
_C\9&)8=F)cF>Z]\L=RH3IS6gaWH40[Y_SOKb=B.Z#(^=&O4JI5,@-AaXJ;L2e@B
A-JXbU5;./X6<=0Sd@SP27geGg?DLSb8=W4V-Jg.^9F(#LUg4g@V<<4SA[A&UK,E
L<:A9eaW<8(gf5(JUXGQY<D\//2^cW&a/Z4E<PFRC&bW=0-bM9U8]bP:+8-CN(6H
&3^Sa-0@3_CY3@F6=U#2/Y?ZSNPETOJ:Y,Ffc@g3ZEf_\?3IW/g#0cMO(H>>O^P?
UW.eM34\0AH[LHAM3C-PQLQePbfg+[dX(.RNc?3[GUL]110P;,900]PaP^:>.JCd
XLacAf2U:,FQY(;QS3G9)K_6DLfR48\3\3W=]D8:M1BfHUD&ME0>YK5[c25d&G\E
0,1;^<(]#fKUG2>>6\&>6CP-GV\]UCA#U/T4.?#TYV\A[Y27F+WMce5141-S\LAN
BJ4#2c=MdTWbXL07)/;_&/:KZ&@;c=2;(FXgITX]QJQdO1_f,DY,H:LZPgHW7bgf
):6<25962]H=JB;/WEJ[=3]5#;O?1NJg\+6+P]JER3XT5KXcD;fU)L#C9f49FA_=
Q1d0EcLH:^B;_:c]Y\&@0[0W<+JN+5]Q/JI#Ye^DY3/K2ReJN&.?UZ]2DdfL#1[V
;[(AL]:4^H<K/4HCE#F^L-6.K-Z9M\)S#?gWa[7G8V9=eG\gR]Ta[F&.<3L?T<SW
I]:+;Y\.26YQ8A/^XP&f.g8WcEH6AVUK+)S2390BebSL&X].D)?IO?]C/SZ(T_E-
DU?YP/&K4^F0/[[VCO#D36^CHTNP3FDOV<V[P#TRG/UW\R)ILWK54PU?geJ9+X^a
ba]QTTg>862LC-LNX\;01BSIX=c-V;VXCf6L=YHY@[?JU;PH_=C.VI82MMS)#S2\
XGT4+Z+B..>&2CCX)2;56H0RM@3D5B:LK\,c.<I>HT@NUWb..+dOL/\Eac>b1_E&
Wg@fS<W_=+H2K1\K?B;JdT],(^Gd--\b>9BT:1E\d8(LV:Q?&</X.H[Fd?^_1/2A
&e--P_dY-d-MTA#_@XZ5&H1a?B(EZeF.dP9TYS,(1V-:d+a&8fP@=:5?77.^ZUWI
<AI+PTHO[LRA.M+c]PY^POYK?958eKT90fV(eA@BIY@E]bM4K[-YC7DE2;#Q(/HM
8X,)Ha:N?VC(;SF1]J,(O@R539a:#(2O,FC\6ET-,O(fS3M]Peg:Xb87bY]@4G?_
31;_fZ1c-<8MUe15EdGV5cOF5_=+b[+13GPYZc\1PeJ]S,;Q>>50I.SHH>NO:61^
d6Le/.BTfQ(U:V1<0eRRPU6\IM])YGbdfE<-0a-d_N66-)=-?YL,1cL+NeQX)P/J
BB86XTX[B__]/L9[fP_7/<EJ[O-IJYY0@W9aL+&Nf690T@OQV^-H,<.2?.\XdF/Y
af;PH9VTI364B\9V#ZP(.KVP>H[:25d4Fd6Q]]MRCXI8XJ8=D]J5BU)_5P<b19d-
&N?\/4b87@ea#OJ3GHc4V#/QQMFH9(DN0.3+8^X6/aBC8,)DL&(GD5ME_]NX<(C?
dM-=M[::XR1=>+IVD&&,Dee?V[^9,@>D\-fF9L/fT.7d/I/>g03U^LHKRV=/67/X
f=5W/Gf+V;X:[/W:X[Z:-.R2PJ?ZUT?2N8bf4X+Gge?8FGEPe)#DYfEegFD+MTOR
)dX#VYO\5ML^-d@/5N;VK.7DI>R1NBJ6Z[Z[9W/=HBEP@40W&IUMdHS)^&f@;US+
6ZZaGd[UFMI;b6&A4N.XZ)@a<GK@:[HRG#[<eaSY((e(G.]JKT5S.MXe^f>RTQ+f
O9e]aFM6Te3UG6e7b.A[=HVda1#d=OE-Wbeb(BDCM7SA:UFAN3LbDIL[FRX#PL4Q
?B+8R.FbUOB&M>gY_E0a_/5b++@7O>IZgV3.3MC,/7JM7WJ\9ZX7)H:M,La54)g>
9^P(+#0I9=,X[ZL878IH&LO&;XQ3+2dH,D0V0eR5IV@(ID+K1:,PNe5#LSUc-@V:
-9XNX8]^LMAeKTT#,/fP4)@,QX4f^K_^6O#Q5F:eH55I38VPAZVF]BJGS6<a]8RD
CLD?c8NMg+KTN;/ZO]3(EH2,Sbd94Q(:]LN?=K((fAJ191cU.X:Y6+RO&\<#Q>/b
ZPeV1Q/@S(c.^.:=dDXAK:DPffO#1S,:=\@@I(7-.(]bO.<?(W;=>UA7X^4I92J,
3aWc:F;GBZDeU+b;7fgD=S&GO,@B44Y7:.+UYQ33cE>XJR[&1@A&+&IFa8bT2YYN
fE[(W]#KOG;>2+_G[0<M<Lf+aN#.HaAYYLSa48[J-YGO]H.gI68DEV,a7W4,4B@4
eU657>LDbZ3f:H##5J+A7ZQ4F/5#4,b+KT^@)9.+e,H3&:62__I(_(O;/SfL/_(R
+F,bWT_Paf#T3#+]E6.YO7><UHNQS2WYd^CgV_X?17OJC8F1DgD5DR^QGHY0:):2
\Z8I>2_O=HK)<RHT^BgB_^^FV-IPS\&64cd/FdD4WOQDY/#ACe9-9+L5Ee2=5+c_
URODZU_Rce8IT6YK\^GHYM3HfX5Xe2B[QfRZ@S>4(OWP9,TY7eWC]c),JN+8N[:W
Z#0;<&:9<LL^Lb(@BN[b/bcU-:<LM21-L;IX/?N6RdDW2LI@6B(A7>?(0f=7(3Hg
<,c/>_KfT5X?#GcKYUE;:M683JM:dcQ;[9;[<GS:ZS0C+QQa4G_ICKYg05G)Y^^V
6UeKe(f1<._NZ(DTP,LE+&8Z<DF=@EQ[c9F61R,B5f:@ENJ34W^cI<KZ5,HUcUG;
>[G#WAU6W6XDLF4X;,2dF,0^O.9a_]OQLR.DA];<CIW_@eB?3S1/Z.1=#X?9R^00
)a2<XLJ002#2@:D7/DV7aGSG7\?L,RDJNef=-[?PX6#+Jdb[;4A[<I,OAg<:+ORY
;]\/[7&->#+#X]:gM8A@cP9g)A<8G1&c\]WBQ&X,)D2]2+SMU9.c\P5eJTM0g6YK
<Hf>Ra4.>_90fF5L,cZdWMd[C>BgS@_[_0C<MOgcb\81JA^LS9YVM+I+1L7#)NKN
6P;7=ac0X0]FdHd&_,3@P^)2^f7N#d/d0B4]^RHc/,LHa@@+,La(-\Qb,4GFW-[9
0DIK5D=RI6aBZ,HeZYELeB1feR4L8gJJK/da(fT8W6>UNFTgE=KLaGcTAE+30=4Q
\&D=ID]QH:eG-:E<NZRBc.6X6\I,O0FP#<HYQ#Ab(])QS5?F-f4]XL;8dc/3VD?f
W1U1-97G-+@Qd@&LC(;LJcQW(S[;6IT4LNc36[3XYNVe<W@9<P3D^\=ODO+0-.bP
I]I_ETd;/L<GS6[P>c>1Bf(WKO/JLEFedbeT],)J@Y.0fOL[:dWXU0L>:O,Xab/S
^^Y+JY:);R:9Zg>7+AB]M8Af2_NS+c<:)1C-6CV_d^_2TPdF)gX\fXH[LVUC,>Q6
3&bT?O49BRNB:#^7BOY+D8[;dL,aB+3=1NJ@^/L+cY+a.]^&A;Z>Pf2+1GPCD[U=
U_DXJDeXEE/]5-(];GYYZfIA?F_/-^PHaWFccI]C-e_VQ2^CGbJ><^c7,E6FU=+O
IP:N&=fP=&[g1>I@.=g4W,<]K.d5KTODe=>#9E#AO+KAV3=[+bEW@14D5+7I6PUB
e8;4P3AA(QLcT50E(N>:_#-YFT>e,+=?&VUD)Da2Rd(NFM39,7L[L]1-<\C?N65S
91ITR?A(V4B(_>#7O_.405aGW(+7ZV\/Q3HZ\MONMFb5Y+]QIT[Y\)fR/9gAeA]?
STU1O@REP+42^_IDMBZ36f_K((4L(eVBX-O@AHB<cg]Y7M6.?C=J_Ig<[EE0[\NO
1O/g4YPK/0I0_BF4]#V0^G)ZYbb69VHD\K67>Y;Y83Nf?O#C;g@(/cEdJUL55+S1
\LFCL@XI1O/Y56>I/:AJ5:L0,,>L@cGCK]1&E@U9W5YJdH<Dg&+GP-UeB09eZIb>
,&bJ.W(cZ8#TOK]-2]VLU<g=BWW^A6F.U?O=S=#Z(:gMGRAG)bR-\:gb1A_<\CL1
N.4QL^83>f+[7J4BYYd6I^BH,]2K4D0()?cO\TRM4?LJ30D>g/<P_8I-G<=Z>Ue@
fE?367ZG1aY.,gWG/IVU#OY_:B.^=,3IAIF+,CEbA4ITY)-[HQ8eI]3Q3;d-3fU#
NGVFT-fd976CK:9((6>-?;&dX6)cLH=2CEV01e,CC6=Y[Q9IAMc,N:VgWS0@A1VP
>NCHZGYC06U:TV4=4>H?>V2gMW=,X].T11YEE-9](OU2A#[.R9-a&ADIWG>Y1IM7
=6RA8V<SRC#Af,T8:MIL\71L]\0H]>)5].CH0#KJd1W-^UA)PD@(R;OYHVc;Q]2L
ZXOP:Ad=a/V1_U9_Sea:S40cU#1)?MWSP=RF;g2RC6T1bAM?#(O;b?V6-NKZRf/?
[985P4dL9RccVYIaZ7PXg9c)gR1)1D_<e@D^F=[\9@E,Y@aV0Fd@Vfd]O-BS+XcM
IHGTT3ACVI>WP-GRFg^?Z3S#)@e:LRX:-[YTJB1X^&Vd^:4U7YXcGKZ//gP/LFd.
@C=g=8fJP_M3JZ#3BH?fD9[S11+CYQ\.&eS6,edf.[1?QbK>K?a&c:+c->4GL&;3
(bTQ1/bX3GWK9MV0:3bS]C-8(OD&.1c#I@gWS+S]Y/M=.9L^?GY9bffE&WZSeFH.
<D(C90/ZJ3;#&B4f6eZ3FW7OY9.LR]<^?1Z#+46c3NDX\\d[C_?DIRgAM#NW>S2[
JIW<+fcUHd.g3M2=R_IWMb?U?X7MM=;:e&CSU3VYLZYAP]93=,^UL\/c4f4Z+]eV
^)f>?=:PMP8EK8c]CSHLHX2\RGZ?eD-AE3.ddG5AFVFM;XEZ,I8Y/8(K;MNPT(ZP
:L0LK([,Kf#e>6Bd<6[TMJgaZ):@abJ3Z-_-;@X#Sgg<1MJ,;+(HEI9_b/B+-O#X
^-b3[;[J3;3:ZA6:,M8@>6C]g+^=[PT)3C_.8dA#e@1@.Z/Hd9a7?38==/JS=^P:
gZ:28^aW@K7gP8-Q::MZ#(gBSK.EPA+Q?3eEE4cG=&&P^gZ0BU5M-Ab=BM8-cV;H
QD_=a]T+dLBd,e^.gP<,BT2d.FLEMSLW=DaIAfJW_b^&gG5,C4C?]TFI3/9_QE&K
XX<R<PXc:#24KDgb@]bU#(IQ2Q>0fgT<,[4FRU34V;Z-RF&.,OO5+61?FF[G+)dL
GXO491ARBX>BgBOg<FSa].bOBNW:/20C10BY/=?+]U9)XM)Z2RIL8+GAC^-?Q=(a
(LU0-VbWSY<]<LcI(aM]gfB<4AeH4E89P/2[/813K=?NdCSf[<e0=(Lf=52<(&GT
)ML3_&]OYa9#QVBOa]2Cf]_H9^J;W25[RR-CMH3PDAE&8>YPP-/YNN&94dIPP>dF
]PaX>@7PJ(M@\N7]_-0NK(CFR4e0EK6M:e\^g/@IAQaCe38LfY:FFN_Y,7eO8Y?a
.SM3NZ,TN]]]Z&=L+TWKBadBK>:Qd3&a,2H)b)(9J@4/8R_SfV9FUPL[.__=B0Xg
./-EK>a;-M7&gZTeG6g169#S4.-;L6..0T@U=A2B:T]([0#)>eX9?OF7])G&>D/g
LZ.3f[W&T]62.UFf\;dFgEJEXPga7?MYgWd<1\(SQFC=OX^a4>5KUAN5^8LcU\0&
\JWTc^NK^7-I^8ZP39acbX&;Q(DI=gBa6B;:-#PXXO0.NaMO),=)#@9LU;G>;:3Q
7F2g5E]9dD2Q<^K#TIGQY69+_8+OWD&/e\gCA\>5+TS&9W[CBEdL+A^_d)3.3D_\
M2::20_3/ZF9I(aGXX5>QWMHKW3]Cc/#25@S+O:;d;b:SfERZO[F]O0(9HVSEV9;
(14;TEPc9g7JS,:2\O\\2\Ug-d7L\CLC<.[,/5c-/##ONK-(QJ+Ta>3;O^#_YFe6
H&UNIV+YU5P5Da5AgP3Ee&a7?\Ka_YTBU.BbYcI7H&D4T[1eA+]^2#CH(_(fTG;J
/AY/CA<\0Q?VET>GV\6X[4XD35bVLON<<\9U34_5e3e9G3S<d#B;>6+_KI#\QX.P
/YQa3@>B4/K-&/fc.8(/Le]GG]@.JL0PCEZO:aY&KKELVaJW@4Z4G.OZ\.PZIa@b
&d>-50MS4DKgKR9g@I\[ZIY\&,#)fO8#VeG;A]bN<.8Z+G>QO(WI(<Kaa+eR=S=Y
.T,O-FL=[5^]3@eS@\ZZ?.JCLI/BbWTdOO2Y=U;?aOfX<?]]ccUSVbRWb^XBFK6S
:0L4bP6<DfEOT+X6ea3eC<+#>)2FRA6Ld5:#N[d+/S\2@>J</Z\Ig:W?>)LP8_^e
GFcOg<3BSF^]cO&/FKK<:W\S1+U1J09F0HSLK87Lg+,GU/S4f0L1.AG@=/0-OAZ>
?DeED:HIM:F:a(gG2(;WNR1Nb9cSBDJb<V7NcA]VAP)00H2:fXJf9(K,@dbbgd.b
bXCVbP2-Z?-dC4?[S;>LFIPfM[F?A8QKK744C5TT-C?0T1Te@:SH[OXG[?8aA(c_
/7+QO(c;P.^JL_4NK,/g[2H>M=M5W:[AG9DKE#H<86X/:(G?,G;R6<RX^dLSBZ]I
S8UK;/;[>0AG<NGJUFG-D_^5K@9WCb2)/O#LFe@P,VJb[0D1Q,?II\UaQHA0.T](
58<4A>XYVOa+TK[PKRJcJcc-\7Yb6,7-SDFBa_NE4gP;&]?bW#bHXK7e7(>?90YW
.29\2Y<.-8\D[-#5\Z>MfU1I[8I^FV1T[<H<77AFOK0\V1c(10bJ#,(.MF9761C9
-50W<bXXWaQ3KEFf=V7LIX6)2,E(Xgb6YPE2d-(fC/+]HM6&H713;-EE<G3S(VKT
:/)2.<>/YA=5A7@gG+1+3)B-UBJS1Bd^e9>\?^<bJX;GZaOaa[NI/DbY5V,f\1[g
BWc]@.P9<E9ZM&4a;PPY=WTS;FRbI6OJD,fXQEeb=./H\)VaA35YTL9^V#a/?W6P
PC5Pc-SUA]4)&,XcX[<HaR9W53X=bO#>(<a(d[LaY)a&ND0Y23S))cJZM>eP=>-b
5XVOK[N&9^0IC4;Rf;.6-N&Z(7XNFOC(Hg0EB8:H7a);PFfD,8V.O^6QH9AX7NFg
@L1QU\E<\KQ](g9EM=BJRc_EV,fB8DSG<=e[N=]=]V?FSRB^8Z:cgR6Yad>OIBfZ
TB.>+<KX@/-&8gH+YUf4\X7)BfHB4#a&[I[QOM507=.G6\aV(9]@:Q@7Qc=A>KAD
5bOE,IJ0EQP+3)WN#Ld7^.P9Y]&:aLBMCeI@_Sa.@W0Y(NVV-Xb7?a0=4ZU?3_?E
AV\?g04O<f=H<\Y=R9]JGM:g>GD0Ie\4-8YJ=15J=]f7JFZ.]S#B7E15(<<5D+2A
5-^/L^(7WIF0//L.O&RFYO^3&U.K=TEb6_\)MIb3I;;<-F6F?^K:QS2/LJbM=Jf9
c:;\@#KR#-E-A(2#P#9:M;ID-gRA&^ZYQ4K1[KLZ/M7I5IA&eO;5]<+]PB46g>Ab
C/Q[GIb_:ZcJ,T:1LE5IUc7@A+AXE[Lb0;=>Me,g_:,-:(d;Y[[W,)E/,Cc6G>NI
ca8eQPGP8(W;e5/LR/JTLd]7ZS^37YJSVbM_@fP2;_0+G^gDK)ab80a6VM8-V5;>
=V;2d/2T7;]6M7>HZ<b4UOH:DJ@8;QUB;(M8TP63,ST=96SHW;BAf;GREQ84,4#_
MSJd02H3;F;LgF&142.&J7Z<@^S_dTcbQ82YVO,8>TWbfb[<0?e4J2P.>:Xfc3,E
:C@T88@C/MYQe59H];2W;cAKO/T+a#9JZf<^Sg+K=XGGOVY:4g;382UbFA(5>X(g
U9XS(.aef#88?/P#eId_>^#Ye_aM^RDQL^:4IC#<2C@CGc01OdR]bbfb/E-A]FV)
=UCR+bAA:-BZHS?Be#@DHGR.@S+HO30+UQG_K+WaN9D#RVMZ/a@I1Q5;V&:72KMY
.,J<U:a7:I93+[gW]/-]Z-UPcg:g\UJSAZ.b=WU,V\dF)e8UQH1bW@9;0gKJ71<2
/#9R;MHe7,;,3HNd#JF6D]>I2-#<c^_57Q+,II=0[#CM<0I@R9X2Te2T.d_IU-3W
&]/NB<f/HIR2T2G]42?=d)9(?WKS_X\9UUKNB>>afSfC<fBQ7SY?#M.&d&IcT8GM
H\:VR.)V_:5e2@JJ^Zg=DOT].769=BC7FP@KP8<G;^T9L^,5+#D#JMHZ+c9X4RTI
d3eHdc43N/BPf23ec_I&4?-Z+UKNUSV.YI+c?c^TVe)(M@B[GC0&-7),RcTdPa,H
R?bN+DTD#X5\4D1VdGNDVSMF9D0MdIKZEQ?PRaE]CV;;8Z3T7Q/].RX4X&]8Y?Zb
H,2<#&HGR0Z=<SL3A)H^(ET3b3_[R03<OC>,A6>^)X<XCG#^<ad6,/eRP,-0-DHM
H5F^=1fI+A_;AgXS<]MHFZC[/5JW7PK6]ZW8aRW..)G\TV/G:@bF;T)/QIEISg&9
MU<]5^:dO=EOfCcbB+3Dd#FWQ=1,K),d,0?_8(Y.1KXMEf<Q1c+6FVdYQ?^#0AcL
Z7g9f0W_7cUIYTYgOIWT1K=>^9;0CYS.4S#B9JK-A)?52:gIWX4XebB-(<LOMc?S
;Z>d;d\XX#1+WFgZH1f[11BD(]g)1Y?D7RYZ2US>J(_#8MCET__P=GYAg/TE#ec]
]fK4eC#D4Y2UVf/@U>TXQ-TO#NW1Pa+(>D>#T=(/_MSW8S:a62/<H4B)J-VSDd=f
SfCXfgLU:5D90\RRZ(MLeEV/SR?-;=MbJC&N31?-&3[P?9IOAF[RG#4-,QD(\dI^
W82,;)Y86P=HK-M)9@IXH,7<<,H/&a/M6JVY,.W@)b^Ne7[>XK/3-Zc]=Jc1S@?3
gGCLJ+Ga23VP)]#aR(W06^^==.60M2Y9dQD.UN^?^dHI6Ad&1T?K@,QgPe7Q9U59
DII,IJBgU+d3Y8N;FQZ;VI\CeJ#d4e,#3gaaAAX9V-YE,^V@6S/>@58W6[@PeLV[
TMd.TUgB05CD:4>Z>1X[++:>)[C@:3A&SGGO#M/,aJVgdOCH#5(Z=M=+/&9A^&)+
M[XD2Sb4^Y>Te5Ab6E3gTH_B+,Jbg=.+8\HX,b:-;N#3I8A4(9fHN#IBO<H/F9Ug
DQT33OgZ/dRIX=P;RO9R;N1=AFO.VS&fE0#.BL&#&c)QHN/1A^7aSY\,R\1PWb^5
-GF&U9IA_(:6-<7(_:IKZ&b[1Da6K=f<855?=GI+[@]54C=HZ8VNA2ba55=:ZZ\/
;6^@TVc-N)00_F+SYTVL/PX5-)SB?UMG:Qe4fHFTdf&1?U-g\g9:N855I1W8&6_>
bY@<5fHH:Mc14ZRF&G[79JGbIVL9X<Z1:I/+bc)4<;N-8QZ#8Z,,HA9T7OD:-W4?
9]9?:&0JO;2Eb1@OZU]fM1@5^5P?3Rb3O^/S2UeE@BD1C+(f)#R@>1g(S0A\?Q0.
X\2^_N<@\K4e9S&NeTB/01W>,Gc\?([TFZ/<74NGO/ZE-ecD5XKX3?X:ZbH2dNd3
(#C.[Q^OH:d.>LI,-R^>O\A^a=8E>JTQ[A(aCMO;Nb_;eQA1A,/g>)O(D?TKMQX&
#D@1.@&X9(;A(J=;CO)R=^g&?TJS-F)?V;LVX<-:ZR<aF7Z.gPcS^BVIc2\#gH:@
C)<@fJ)F::>4/#6/A+IU&J_De(4,919/eD:H&d68G(Y@[A;B<,[K=^4O1NY#=8c@
U:/0fbH4WDab6&=+[aK=50D4?Yag;AMd7a;2DLP=1Ng<;?8KRRJ5[IW5)Tb^H@4S
]4K3OQ_)7&6>LN+,\4IU3cHa0g^:((I=G/_XKVG=B,<[TMW7O1M]f,,7d,A&(2+P
A?\O)KI3[E2fM:^S/7+Ed:c(]Uf99\3W^7)TM[@R5,,HQS&-g]EKOWD\JZa[,/_(
;J62M,?E&]C;-b\F/[3=#QFHe\OPV^g&SVX4YQ[<A>3_Yb#a&H=B-L_.CU2^e7QT
=JbM23(P^4FN/&-,H5^XT2-APQ,:N&U@B,78W#[B:a:8>)JVcBe\3g/><:aV500+
ZX/9K.<a-3gCWNL\7#a2FceI@HY5b&f>Y?R6:OFD2U2UW3TcO<#OHaD\F5(cX.0H
K;I]@:EJ^OZ.YZDb459-6IY@5VBc73#2/9<bI(&FPbBf)_FUY._F4+N1beZ2,/2Y
B2aA:0>(O(EcB2.>#SGNAFFQ/D+Q7\-<A@9+BCOVeaK:KZ7g99RJ1fN>TDaWfL?I
@M5KgD_]X4B^3GO=5:c-6=f_Q:)I<L3HK,QGA/P<0_0SU4=F@&MPed;>eWefM8D?
IJ<N3YM<L0Z\Y9AG^ac5TLf+V;>6_ZX]7e.)I2-9eN+[1g@<a5&ccE@\bG2#1(VY
SKAT(ZGCL+&6N7_AU5LC^+.YK^6O5L8[1BA/V\db-5N2/^f7=-J4FNK>5eI[Vb)3
.;@A@58(C9H/J#Q7BES/5[;dT9(()LJRHG@fOHGNc4S&R/M(A-#bD6Y>dK@b;NE.
JMO=4We(#gPE)F2gf9(:T[M1[Ac>R7(E@?a#aN#S4-?FG]P/LQ,P.KO5=.D)0D?<
bB6Pbb;f<+G#_UMRW;#67CQBdP8\VCHQV:U0(feTaFFL8b8.O.&7G+KK=\8V/S)P
1Y2e2=/A&8R2H\F2L37@Xb&Wc0ELFSKPIYO=39Y4Afg_[Q]V06FX4AM3)1gfZ1DH
2XS1/8B;MWLBIMU8O6TBHQ<P2_UD[cYG6bW\EOf;P4NQd)@LO?@5Y?XB+?:8T4O)
g8Afg0@\Q5Ne4<K<BP;^;T^:P2.D_,0,AI3DaQM3X-\QUCE_b_GMg6C&XNTJG]f=
GHPf#dLGg1R<f5SG_ZO]+[3?]Le=AfK&BG<:bBf8]4?:bc9(e6^Qb;b&+S<DQA5W
eOL.JI=SR.S->EFbSR>ZU+O5c1eI2#=2FID/6DID_4-0e/:a(4/YPeAL96X-.RU5
;0:.H<N(ad4(TdAV^]+.<e0G2;PLbdB]#3egG?W,4dEGLTKHPYL.D0F<X0HWK\CF
Y1O5<I>61U6A_R5M=aT;XNca>(2=g&I25TW9@4^=^?&E&D<&)QA&^N]0_P]+(fM_
-b)HLS1_&N#GSAZ53XFQ/[,XR>f.31F#3G,(1D>=1;]8-6SaL(.gR^<01#VMSaS+
aCY)VOMbI6@1@(HB34(RKHN2&+U)L8V;8Te_2>T]TC@a^U>Ye3RB9D+Z,K8cSXPL
d/^-EaCZGOUO3[g5U4@6G>PD,e-KQ/ZHP_Q+TR-P[P8^f6-Q1=>;fgNID+O+KJ(f
T:P/EIM5P,,I/eC3e1:aRUVcE[VL-2X7E=&a0\&bSfgYa7Q4^.-86Bb[Hf(G.d]E
6EL=R;H<TJH\QUPE)^_NE:_AFS[CIY9SW\\VOaE&We/QKAP4DV;14&F=BF65,>S+
-^357FG4V?]7^KSS>SEWbeXN)^X_WOed+X^JK?#OeLL/70gSF<Lb,JbS7ed(_#X#
V/&d2V9cBCM)YF039f6b#-AT:dDKGK-45(N(&S)90;6GgA>.:)@EA@&]0DW/Q97^
Bd^ZUgQcQG-I@bQ+]>SF7GbH4]N(D=YC[=5FSL2d[/>/7B&UD?S:..C_QgQT<H>U
&7BSOV3:6WaQd8#=B37MZS;R#edS.?X7POKZK+@JG1,DQg[D=T?;0;==0>8UcRB2
I585?@_OA2Q;1-4,2[gWT^eUMNM>(2D46?A-]K;O6_Xc65fP#HVcc,0L<R4,6PPN
d<,1XV0H9a95KG+.C_#9_Bg+e.]b[+bQ._ZY6=e@Lc-7\+6F:Z)J]P>>aY1FMRED
ST<M#6@6QL2#1S?<4[/8+YLG;VJ419a/>d0#R0,5P&YCZ&[/W095AgZ(+S74_gX1
e7=R-VY]]\e/Y[,U64Xd#\]Y&2^Yb4PKEc,C\7?3T:8I0WW;XMXGL#::Nd;Pb\4K
:(LGdYW&ZW8OP>F(/#DZX/RC>O1Y<25aFD7=>SR1fC;=1#LDLQ9(A=4d+?@87GJ]
MR0bLE+4\a>@e++d(OJEB^:^GE3BJF>f1S?V5#LAa&)#+#621Q.RD(C?DL=OAIbQ
4MZ9:g:,K?0OQ._)BTNY[<OY3e9BeJ<R@/4QVHK^UTRa-JDL<1HRP/GGaY4R]629
\4.?(^1.8#RKF?I;]X&H;+67@-Q)C[</;>:(3:]d6?beI<_QCY](4CF1E>]SF2G&
G5W)&34Y-ea]H?fRB1X(H]e+c&1&[5=WH1=CJB\(D/_(gO^7&<ZBC9,42GBJL6BH
=E2E\AM\Ca^J4\^Q8Pe)dDKY#CP4.Y]fe4R93_CT.K;a7=S0NR;SE7(T3-[)H@Hg
^(FS>BI^_gbM-RQ;2:+SZ2/4ZXUSP:A73@\^A8HM<-BB6>1F9FH)799L^A>UG3V\
^X8Z=#M,gAL=cAIM/&8SNJA<00N8cP8d=U1^P+QN5,>NQ_5,LCec^488-UQVQ3fP
3=Q+RF-E<XJZ66D?]ZVg1D\\G;0DT:O7.9B,b\.)IYEONA5XdI?._N(GDF/K4(<7
GJ_V;P\^d+/49X2Yf6Wac#2292C2A_]A3\^YU;/6<(\@6&>F<R]2)/VYO4_-,@0X
NW?/[.CIHJ:\[QPJV]d6(\-DZ+A<Rb\^?UBN=[C635[Aa+FF:51<\UA3=0->gGGG
OX0T+KAP<82eQf/)EcEC&^NX,210#+R-&b\XCFVEPd?W7fQGTALERKIU25K(ZaNb
f+:TG:bF@2H1^ISUbSYVA(]3b,B?1JYH0D@KWS5UUVSW-^e;RH2XGbF@eAQ\L7_a
[Y(b/6Q+ZB\-(&2HA59f0HD90DgINFLN<VEH5(gBUX4c:>)2L3)=Lf<:A_+^51-e
>M7XdX97040_:=/_SN&7L6RW=TbgC[fNf,AFg?35JZM&J3W]d@/;b5Te\f@beJ6g
/BS+S=MFGA8YB4VAJ/I2:0fbD2P:9)?DEV?<^FGV+C\d4:dAG36FKOfZQJ=;KaQQ
4<U:##3QENS/#R_&b8O^XbfHN(;B+,+<?JaIG;NK1,QXE,8(>PYZ/J:M6-Y/=2F#
=&:?JfQb]<]1A]#M[41Ia=6-^FbD#<7S7E&(7ZT(M2]e0/6LBS[T6Db&GZ942JcD
03A/F2CDAG^c(<_d+VR55+SX6b9.fSAE0Y(KT@O-d;+K_\7Z5#Cg:I&HA_1NbIU&
83,.cNXM;,DeL]aY:RbQTD9&2C05VN3W_\@0EX4])0GMeJbJBD,0aP.g.JQLWYAa
^M)_<aXIPG5X(N(8CUYR\GRaYWAV=&@dV?GS#TPXG25/B.2QI^DKb5@YHJAJ?S6(
Qe&B(@LY0UV^AC:CFPNgO]F\J?XD&E4HPRe3;bgcA&;R9=Uf)VO<E&.X/;6Q^FM:
,8--DO7)a\b)5d29<e(^R6LO-\gHZ5f[/2/^\/.&S90.X?Ae[WC-a#PQ(RQTK];g
Z]#;\e^c0;;/XCEc6d3VM9Q,3;f]/QHPX^@]<KP5a1D<9T<<^4-eQ:RH:Z+#(ce2
UMK5IZ^)N8ec4<(g[0PE4+:93;gK[X6,TL;UG^&B#GHR+8KJ^B;JS7eU#:YP#/,I
Z3[QLP(Xg9U,[UFY(Ud&a;GI2OY>GbVJ;/;8/a4?+\UZEM]0(U6ac?2V9-[c<Zc=
D^;U>b-O^<]YRW=(eW5[N#^dX@MY[,ZH_]e;E:0)I@?;f.T]NcWHHM83:<D;7X,a
T.-,dS(cO?Y:7V)BgT6]07J&\-g#.6P&>XeG;G.+(>36Z9+ZB3H?0?b?=E\8=.4O
L4IbHRbXE25^e:APQ=Pd-K,4[K@AW[+0KJ+g)^Q7^<Z3D9PV-c7ZNd2VAHHCKR&_
44bUG4dJg-6OTQT4SI]fA2T:<-=EYUD>8a]2O_@^,;B<M<.b&2+O:ef-ZXB<Q;.G
Y<cO<K;Y^S4=ITJO80Z)0PUR_+FY0Z1D/f60B_0<R;2fT6AR<F&RHbRbA5<=<Gbf
B6@6,&/7.f:^@0H\H&M8;1E-\-KU>?:U#;&E>GVcQC@aA868)Eb5ge6W7NQcZWUX
W)-UaNWP_aF9P8/GD1XD&L#[:U67N#B/B@A8X>J/)-[-:F,Z;ER+a=>#KM2&-fW3
ES1b&W8+:-SAW^)e>ZSg,&CBQTX#=VYc59IDX>BOdX?Xb]11&X0E>\;G^3,YP0P1
Adf&74fLa-LZF5H[B<P/S8](UB#N.:G8WY^gFLR&0-ZD3SKZKV9:7OD5AO?)M3JA
42Vf8b]LVH4H-4#(B,FSGc89NObV6)=W,3\SF/_(?36BM<@#fIW;662KSUe0Gd8K
&NKT7_L@F&CE\cW?SJK0Ea=L6?4D;EI@FX#_-H88e:I.E<:d(U#SDcg]g@Sdcce)
cN&>G/8HJ^/Jd(H1IbB7d?Ff[aO0V6C1/I--d9[dVO<;_E7]T]QK;=885:E=<S\g
),U^K\<R,6PR\IME_3:#fSRD5UYN.]4>U-K&T-J\?#edM]CGd\O>,dLPG8U5C-YT
5Z2BfGFFB^E2,.c.73(OAR?<@<>V7))A^fOVd8eGWUX5c8MR\:>,eAGUD@#S2M:3
Zd;;@ABQc_?;6a=3a<+(Gb##H,QF6:&>7f9TYJa7^=6EZ@#4\(R9>(7&?]CA?aOe
Ua#P=]0+,V?eX&KBF\0d8,:YP9&dZ1Z0fJDKO=W(W^<6W<9/1WH4_1;,JQ;@YMA,
/T:]0,c91EDE\fEV:G9gJL5E#>E_?U)8&&JPeJDZI0@-(f4^G6/AAE=VV^KUeea&
&1ZU3Sc2>B0+D&3PM31CDNN>JS;,beBAH2@PNHDGTEAT2N4N>^>(_bDPde9)_F=]
<dC2(5<M(cMgPI?[N8d;Y[5<Q4R4CM_^SeSAW)[(S/=.?JO55[2D7HDJ>I#==>-1
Z?DB1-g]&4C7DUA7Y]d>_.D)2_PD2D(_-+&[C#V0.2dWUc#Yb&S4a#c]ZRJ?69XA
L-UR5Vc6g((ZS0I)9db1NO>RdR+3]E7@.:9=ES[OFD+:->W(>(WZGTRGXCHGIUEB
-bbP,d9;-&P0^9GMTL;(=A-N\JX>(a5b6eEVUI(B=f;d5XTC1H+RC#[c@214aK-=
_A]KDMFYFCY\)eS\BU9:GF1>L:,58A@56F+J05\C>_5OSB-XR&I#F78GIZ5P?LU,
O=.7(YcQ@SNLUAEda2X6S8;3TH(&EGR,EbZU#=4\R>JFT#:>@(=fg-dAGDDL4A_[
Q86@8U;BgN6O]>>N(0G1BO-DLMc81KK2Ze;P0(WW&+02@3UXFgbe8^Z90/fH0Gf:
[;<B#GE3Q/CMWaF8@U>X)&+d^K)98YH9>S]68D2S_,49>_?-&Z-S/F<FY\</^c-Y
8e25Q/#,aN,OSacdATdPeXa^=N<S@:YX.1F0/B&HQb.V^YMQM5SP..4P&-VK#S93
IOfW6Q3CE4ICD(BJ:,aJDF_(Vg>A&SMRL)Kd\FFcQ\KcYI4Zg8<\2C6HL889A,0B
N\-QHUU_.&Gf(<BaD/P0R,SEWHH>L]:72.H73P:6+>b]@<cP.=1=Qe_FN8^P?.PB
]Wf3;4)Pe2U->=ZXV0E:&>AT8,N<F@N@01_-)5-YN5df6YB\<UXCR^?AD>B5D^Qc
T;a(=(&7-+aT&VYN;U=Sc0R[[5dYS;DcCKCD++eQ&,DRf[R7J6SbHG,X)>WJK9gO
#=P,C27_?R_B-U:WP7fc]PNHbDc0]XaL+:7/9<)1f#VV<PN.eOK_,KZX,gdK@0GS
ddW/OH7Z^MJJ@[ES:@=2:+=&\PVZ\UU5d95SZ9>?/J]9/Z-P[gFd2W&\MaX6W,)[
SK68G;0UOHF=WO_2;[M)D7)#@3-&B1<FR?;+&4DSBH2A<S0Fe-CPg\_+?cD/f2)W
b5<T_]<TN[4B]F.HcJ&bHS6TAc@gS;RBfXbER2+)1;[3(G\Y<PX6&d:eSL/,V5_d
ACY#UW@Gb./H=J]93&:[&KJ8KB].HT:,G[,f7.^9CXJ(]-5,XZF</GL[6Bb@U)M&
gdDfcD0SaJ@QB2T+9\2N7LNX7R27I\R^U/-/P)Dd)>:#9f#U&CgbVP:)C\Fg(UV0
f5U;>@gMaGXa69;OI(f+TFeYba59OG[U.M>[OCIOHS.Y+S]>B]0=.>g^R;7cIg91
JFa;)>:?96d2Eb:Bb+6>Yb4+C>9))4FeWY5S^6W>,E-GEC:Z?DQU:5gHe@_Q4&d2
0M\=[KOT872[X98C0g,?f(FW3\U(&3Q7Q4-_Q#.9Z=?X&,7.0--K0f/I?K;4WbHL
/Z?]081a\;WXKf&f\3AGS^N9MM)?TdXWcX]^#O-1FV>_<I;Zfg0bO+@Megde^cVI
@E^7c:M,.M9NAQXg&9PS-[-4[N#LF8M__dV)@KDJEB3<(,[A_eIa]2T<a;J283+e
RZ=)2Z9?UY27KKEN@)I)AJ&]66#QYN@W-2IGfCHJO?H03+6Q@=\?(2/W-M5Ef^GM
Q(gaC.S>,-27>BO>B[_O-TS;Q.IU.@[Ue.gU;Gg<baB[HVT^9MeABXU3BJD:L4MU
S5,5=5&fE\D.>;f-RA9+#g3WCIOJgR94(P@Rf8:F[+:A91Q>@0DX23Rf(O1RD\0X
DZ4I3M0d.2U1<N&VU+D2_-OEFS1b&_R1UUg#7G4L;KLJaeV^+MBGGA7#Jd=(8Y61
8)--6;^GeM:XcK?77GNY_CXXD(8+Xf>OQ#:GE[E5g2JY_OLGP>CVXUd)f0&>?Q;?
W8K/6S^4bOM#I#-GEc(AT?]5AbR3X&7\TK(d[)UI[3Zg09;QX9WL3fMZOW1eDT:#
SWVGM&=YG25beS;1?&33CUQT^A;1IL+I+8060C#4=_b)72GKYLB?G=G=4]B^d-@Q
Z_IHD_N7W?LPO9\8X9dA)&.KI\B.._\8+:gVN2^:=M\.cCD?-J)5e[(,JKJU,fGV
]./g;P[B<.2;&;MI&_N7\S-7e[Y_c[5&AgI^,MH8-L(b82AF)030EJ_^<W&R6ZB:
3H\-aG##YT.H]TXOOI-;6(5E^QO]N(0T\)LY]YZKG9#>P2OfP#>+K-#:DZ=RQ1ZZ
4.U-WMa-:(#]BMJB>=DgW[4=&cQ;_aZ,060f:3fE&b2)CA^9b8O<19b2=3=LX==I
Wc@@;?:=ZCU2JX=WaP0WU=QI#N?I66I#/#8[<fX5BWE&59c:A\0E.Q8=D;WAbeHa
L(M]X796Hf)M_X<e6S668g\gSTRGW4OQ0Ge6OR&D@ZEN=dT;86(X2LMC_BdM+1-+
Za\gRCO9TZ3X&WfC8WZc9S5dXHe@)(.6S_\N:?DU9aQa[BD[MG<ScYd.YCE))6OJ
0T[(X<V8ZeC^2\+.2R5@(E;4BX.SX3[=aU(A>JU:+EM=1/95,1&9^dB)5E8R:b<N
PHM0c-RRb6?Ae9g>,[VRZeR>c=&<e8Q(ZP=DO[dIN>QYb(G9ATcc/-W1/>WNJLIQ
7FeP\(28AL1gS\fQ#a[M-d^IU(,:B[?E:&(:&>V5XMf^B]Cgf#4D:FdVV&MKeJ2&
=O\fQ1O.9EG_1R.PfCL8G^LBHUWI(4(;gC,[77J]\e>g9_c(62J2L[C/O)26>^:=
SagFLUVT9[_NCXCG3Y#S0&^O/ARVL.@OU.c7T)N6L673U1-b=HNLb,fE:KA8Ig=b
K/\FDbfe&^X_ZaACKDBIa,eaE@<Z=VENU(d0d0#Ka0>W7C7[^GQ)#UD7\KEE3SOW
H29L1+e/U>cJ9Xb8V4<;VbS+/XY6=c/7_#_(DV]gfJ?,]dRP#J2Pa.P):R5e<)#&
&^MINS;R;#_)@70VT8)3gg,NEfO\^B8>MR;2eV>V-0UA8U:1\YY7g)5g>>/W+-II
HQ?T=aCDaa+IL:E?W&_cBW4H^6U>,@:U8YUDBQ-;dYAUaBEP^BS@8CKFS/fF1V/M
gM(cY=&PEFR2b?KIgPM./N[J<J9TI,DdW1Q^Zb]=;[BG38eH;FP6_e<+GH94TIc9
?GHPSUeQ:F_RB><?Gg)OdNIBY/YT31\bP<Dg-P<.F&#>AK3gSaJ/g4K6H6UR1V<A
5cQ?6IZC143;Y6>9^QT?8<?<^.;S_32cELAUg4Tb<7(fS=CH79/L)<&7?UD^9V>R
9?4<feHR-H-X0+S8Y_9G/KB7C+/4^2N<41429N@6BKeTeYZ1LGdZ2XR)VGYX1FNS
SM2:(61T(E=VR/\^,,HVT1=LY_,</F5(?Jc.aDCA&B)O3A++<4P-]b&TLX,3@+TV
T5X<7TL6P_S=[@D/DRGE1(;Q3G5D]3]]/&Ue,TXd9XL)VIGc\c:(_V:0e0]IR++a
f1\##bG&[N9EX5AH6X7B.H>B@R1,L6/+P4cQQV;=FH=DRAK58D#PAY[-XMSFIO7+
aH_L]GTA3AA3QQV(GECQUOb^Y3)?eDe-Z&<)AVJ)^QJRZcJdS0DGKY?#/3Y+aRI_
(MJL9WBP85Zf3a1MUEHdGf+[XW<7UTU5WFe3JJ<E)MK7G+-EC=G6:#K=NDEM,]a<
UK.aF\:H53e_KgS;fc7_<(^P[6,cf0e<>-eT7QXC<>F^DKRYYL^9;A0:MI-^J[Aa
<0HJLI1JD^0VZCRA-Kd/03LP1.K]O-#aWcCXA\2T9E:AR-gFSCg)Pfc_>2]A\0B8
(g\2eBVDBJeg:^,^E+Y5#=3TMSgXLgO<9HKfGWFSW(<B.[ecedK7+Ae6#0bS9PN0
OS&Hf3JWMbQgYC-[6NfZ&YV7].]TZ,=d3(UB5QV\e3OFQ;F5J6fKSJ8.+TO\HLJ-
cPf)@AH.^aaAG9(2P^=&:RXP0DWc6VPba;b\<,^R(#dJ=ADD#E9RgSKGQS])<Qa^
UWcF\cY?VBV#ZU8#QL,8/bUAE>RK?Q5/IVDJ0\W;ZS7VOLf0G1R2e#_8a?<OH#Nd
EIE]G.C=#9d9,GBW5[@P3gbB6L;]X<DWe,SL4:aCO7W1>Z8A[Y0)]NDYRX]/f8WP
S\fX(ZO8P5QBN(VN)Ra6:<WB:F+SR#F<VI&0A,)\V:^+VDXNB6H59G.GS5:D_6^D
#bT6G(F]SJ1Lb8[.04?B/TZL8N-SH9PLX(:,,^R0.gUYWV3Z+#.,F&[GEIH;D5dY
:0MA\eE.>T0<[=N=]4,<8?/^\81fdV@]FAGGE9]JSb,<E)+_I0ReB&Dgg9eY&8ZV
UTRJ<b_PG[=MK5?M9HUNB9Tc9\/bRePLP&.,dO_O,gP=I8.9eJR9J+)=QE4YNE(b
NVOOgRV;AAOCRffY&PB;^c<M-c(0;97gJJ0IN;L+WM@OA>^:I0R7+-<<\KOe=9_B
cJKCa-g&<D0M9W(Z(>3PNCT[f5^<YP48dcQfM\8EWB6A<04KgD3QNZTE,,eZ=Fa:
eF\<T-[TL\QR)H(T@aWQOgP_V<99B;8HP8fg1-R7)RJ-8AbUX)V;/?,Zd\9+XZNV
eD<&WHcP=^MfeF&1]@-&#J0\&9I3=&B5,:P637:A&Q0Paged5J==c/[O;]b=FcB5
ec-AD9=(HY#7TFQR8C_CV@3#f]7@>a&/[ba)/X-^2b;_5SYB]<Q(6W(33-J>XcDV
:_;Q68=/ZUM=a4R0A;K;2(,-KegM.P_H3NZJ<MHQN-,P+91G]Qd_B5>N@[>aecZH
3+,&8#.<XDT)S.P\/FaZ65X7O,[f2B5QIU6IGWZ5eb^^+3I87(Id8]dT?R?81JUA
2ab0E,Z3b6fH]ET0G4@.<^,13cfIK1^ZeZW8304eBL_RZ\;6_QggA_8J32&XRVP9
fGPC:Vc(\9[&Y\826O->7[Q29X</VQ&P+3d/?/3=We3I2D1K@3GM?F,f7(^U&SSR
b+6C(SYO3[UM@Y)dfW(I=O<g2]4H(b(/3RZ@&27aS>RCU_^2A^d(^aZ2KCW0EH21
H@45+PD\@c43]RU912eH,\L@TWXVOD8-:MNP2#I/b49/_9@\)BUHC>1=M+[2Ub)5
a0-7EgeAOK4?dT<Oa6OZUK(A/-^aF>5>e)Sa)?;9IgC=C@JOT6Hg@V:Q,M3[6]He
AR)KA115NUBA]P=7C5/KXDKVWMOJ\\WL_M)/Q&HeJ07CT@KV6W&Z\LUdfNRQO?]B
_Q=LCS;;4[9U1@/L4\H)USf3c\_KDZ0B@d6?>LS7R)-7)VO>E,KEC;;a1BdB8(CF
48Q0)M[TLST9&4e0#;;KC:Q6<CEA?W^BGc=B,^1_a@AP=B0UEfNN90c>X:1-4/Mg
P)37;gCH-<A9;_>XPd,eLR^-4d,XTcgScd#A+RW3d>Y&d8[Pa(9&9UV0,E22HUV6
<^GVD>3T.68BV-=ODGM=:9:\N;F9a_(Q)A2U.D2EHCf1(.7XYbYf2VKCE(c^C^e-
#a9f.=6T;>(AJa95e89&,]5;,gQJ8W/0b=@aBMZEUV^.H#4?4XW:6dKG_L(P+Y;(
eMK?U)f=_NB=1MLH70+e]\e.00DfC&]b8MMgH,L0ZV^S8UTZ9]5@D>/#[75X1MIR
+3>/61_UN::ZN5E1#I7L(d+ZC+]cB;+eWCE@e^G>cgI6A,c+].,d9RE/fGP?g?aU
C1#27XCKSeR&I07-19TCc1A-V4=abS7,;=SJ7;_D7(D-7UFAbT+Ug?<&E9O[.SAg
-W,@E#><^fb;S+K,fD4J\5b:eB[(1U7C]1(e9_g[JZT3/=?<8#9:P<P9RdT_OcN8
Af;Y[RFPE;7D>T4+//]d(\1CIM=Q(YH?V-7PE47.Y;LV/.7Y[bY3Q?WZ@VP9R49.
=&T_9C>I<VQ/<R,M.S_V7_.HM3(2#L#=)gHF51][ZeY;5AgH&Y/?:WGaYfI@fP8E
;,4Z19X5:>\<VWO\6()R7_CLWaG<6e,^A0H62^OBL?<?a+:^6/:;&RK2S4UF<-Vb
#]UBbD5E:1[5cbEVSbd[.G+aZ16(H-YBf88&#Y^S/LH/f,N>_G/Ea9Aa.EZM,]c+
e6OC^9?D)VV?9A,AIT>[R7V?26)]=MMY>IeMP+NgPbPXFF#IU[CM^GAN,@PQ,;_J
)P)HQT2:#+RH0O,D&\VGRgW3_BCa93A5;ML48HGdZV=,X2_Q6?V^8>/KeEVggGMY
>ddGMS\]&RG&0(c=(I^3M+/9-DJXJR&.RdeTKa#LCZ7?Y)6ZZGGBd;g3U@QA:NYV
+VLA0cDf^M.WPK4\#)cY\6L@VG@a[gCHXcTN58H6Q/^S7ea.LgAbKg]a<1[J-A96
RL:eH-)PAJ-.dJ.c69R6K@_fGL?S=J,Xa:0IaOD]_WdF&5X\]IC,XNGZ7PKS>;R^
e?>6,+L0IQ#X\I4IWIYaC^@AR]@&&G46C//KN7BUK]bMI_eRgJQfFXZP)TRd2#F@
#1N_Q=3J:IV](LMT?W.0N.>=SYU1g0:F:;c09b9+T2gE#((F;=O(U[OYUc9gX5Db
P4S(JR@F5g.\4b(94-Y2U0284#CPO6ce<EK[WF+C+8JV;4EOM6bRH0dNL5>&&L3@
)VBK^9AMgPVV5&-OU;[\CRVgDdM(IRIM4[_WT3bU[Xc52#SG+D\>OJTKT5Z0c(U4
UFS:VP)-fH5C;OdEfYNF65[5aX-HQ&&:?+Ob5EB1?+e.fU6TTAN\OI:]4T?7;GEP
ZOF0R9CGKBB2;c7L?NTcY\TE(7U=fSPB->=[cEKZ(PfMJL6;3#Hg-f-B_Jf(C\WX
g_-g-IX(d7K;b<_#OF<aKF+FCa;92#Y9\[b\DGC/7Q6#J>5BbgU:^00:9&;939E5
7AQNPQR<.e0aG/KM0]<:1/H99_f6c_2_gQXPLNfY847P+Y^&^)U-V[\8/9V1HJ##
SJ/AgaO6UYVT+H+4aY2,Cb&IHg.K2CEc(eF/+)EY=fUO=Sf,AgMII&e;a;.B\gDE
3M+AE)/3WHYN]#Z0;_./,/NEF^N)R9X#PU23[DCfA;^ACMA/?c6430@@D[Y7dCIR
g3d/K<4^7P,(6;^/896SOX6TfUR@H&af[[,Z/T2Z+Y#YV&X1#E#<F<<Rb3SOD@,:
e8L:3+9I]C^cA?M[8VGMQ&0+^I#9fJLGOPO6Z[U,Sec.C&3K)<;:-\(EaG_&BKXP
&dX2)P>_[1U?M;^X?Q@;b)1;,STd^)^?8B^F7SD(5B=_Y]>c1XI4Y/WS](6SSVFL
_27UB)F<FN9ZcHD4EJ:[e@CVIUYE@[cM[Q(0fMa1FQADg&7/bBQ(QWZ(2PBI?33C
5/KJe1/SgeP8,Wd/.Q>9Q-b=]T[(1V,O?;+DfD2S,7L)<07ET3a5D;I:/@4P/[T=
CdIZD5I6&,]V7T:UfXOSI>g>Y:&YTQ3]_4T.\<+4?2_5D2\Y0\GeS2L?GcV>fY@4
)Q>&T#,T5<,HfdNd+b\#^>E[=gbd0&@(;LZ7UTX1dQgMa/D+RR-/cDCGD&R7Y3T3
g5^e[-KKBf2>4gRe<GI(PPO7^fFZ?^VJD\K-\;JZe9a)cZcAE+^(T,KQD@^[@GED
X1A\B3dM.QIA(.M#e(MT2M8e,TcQ-d)Pc2PcIa+GS&6MNaW.Z12g,)\;N+QIUdcc
LAaWIF6eeA?J:-8)H]JW//#_,(R,0)Zc)QKY3:9VX<_X;FLMKK^872LP&[^U45#C
?6&5-+,^)C]TQaM7\X&8[[NMJNg2dZ-<3Z>Cc:MCLFA;?)\+7g15N;O&CNe,Pf:1
BH-FO5J831-d-P60U,Q9gR[fNT/9GP]2H9BM&3e&T.98AeY+0HRH2;eLL]@:e444
QY3FPLcN:KD4bEFQ:=N8be#HJ1::,C[c-[<4:EW&KMf#1L5(QXGWd#?OBP-D5RPQ
I8\#DJ,@>d[@C]JLY1KT^]I@C2^O]AOTK\Re\N9gL-,^U<5JH5?C#W\B1;3=g>>7
Y^4fYBeV5V4=\&7/#17ZgeGFPMIFK).R?4e<UE32N7LQ-P[a#C<>d]IZ@^\Z2(/6
J-d#<SGHQ.2:=:.?M>4g;&],2:+SXRD?<a3UEV]<#U.13-OBHc:\)c9,UTLB8)<1
D;E#4_L61P(eLDB8]R&O/aeK8FL_^--7X@\:+\/,SbZK?.=g79^f:K[>VNO@&S1]
ONA)T0B50?,^E>][e,QDZI?d<>Df#D7KG(YWBF7W_/4;>dTaT?c9?&2_2G2VIA&S
W[>g4b720<?GO^2VaAXZS22P0b(^=XE,Y9]DDf4V_12A96gd\&DQ5]-;(f&)UQKI
7GEeFB2LY>42UXK8BH11(?-^)3Y_[XfeJB\g)@I),ff@#a_:<fBV_7:Y=WCYN165
;L?b@#33C=Z[c<?JKc.g]39+QGZ25:VUY]\[OJX&6>JAc)4\)24S?HF@1QO?(W]D
TAKc4NP[WEO#IE@;/>fM14]E;gaGbG2aa+c\aWFSR/N+SPK-W)SMKfOH7<_PRQ0Q
5b;5U2;-,?(/Gg(b3=>6?&=/N:@c;3>E6;7f;PF;PEX(3GXQ=Q=&PX^9_21:Y=9Q
HZXM>/\O4;HGdHR1M+S+0RY=1M(4d2bNaDMLFTU?09O2ZTGHdV&2U@;=+@OZ5N:(
=Q<(+Z1g:,d.<B#5EA(2:d4bV-2GDg.1YURB/1S55SZ@[67P)9?_CM?6gIUUTg-.
JAc=:@QMaUM80=/>(4P4bLNGS_N4a0P23(Uc()ERNNFXRgVAK=.;9E@LW/R&aI5&
Yc0_;316d<4C@;U+(2-d:FYbCN2Gd4(HHZ?24.6M7ASL[3d+=,S/6=.0&ZWO?JD(
:JY:WKScJAEI)7Q2W9;T9C1-RN>(OdX-ScH>dXY3JefZ:Q(/^C6bG69L.D+ddRQU
c#V^UIM-J:<P&<WOV;118Kaa45gbS5dBE/:aNb8&1IE1MDNY)JM1R2CY?3F&?G<:
X;#:V43C;f\VWJXZAe5<&^c[^L\^VN?FOS6@H<->=PbHV4g-ae)6NXIN[;,SOL[Q
A^JOR#AW[Nc?H6S:c6.Z-;g;S.NIC,_9eSGe5V,E[F<R-d2>Ud+Y:3Q8;GL3Z22]
R[ROfUGM>K7;T7I7ZHQ-c&C?[3NK>Ce6S(\SAeK:83DD<NK_3>&KTN:>,d?E-SIA
=B/7g?4I.b5#DK+;E<=,H<eZ-;LNWG(LL<f0ABI1_(;3f\##Q6F5c+9N<(X0YSB\
Y3_A0:T\AS.2AY]EQGA:cJ^gV;YW>F>00PKD2L876?0Ub>0.YbBFULYg:7097@4_
>WGQe;O60Z&I7]8>F/eDH6UGG)VBD5@R7]g0>a3RLf@3>BO;V>f^55:UFI-A4^(+
H>TTQ,aHcSW+<N_1FB,E?YdDBAQO(QBB2]GD@NE:7+UI8GTc6c;DJF(C[,b+2//^
/GaTg^I2@#UeeR\6f&I31+#]/bJ_I,<F_UTNHXUbg8&S:4(g()HY/.MJ/eLH#6E>
Kgb+cWZGG^1FG41?bf;G]MYZ0:)RM\R@/IX?f3+#&GPLYQ.gZ0<3&W.gJC>X9M>[
S-6>XE;NI/DT5&<=_5[/BDDOK=[RTY2033K1:ZQXOSA&AeVH7\;@QcK5/J5U?Z=K
(R9@==C9f=N23HR3<@-?cFEQ+dQ1YR,46?+)V>TVTV,R:Z^NFZ9Y<5+F5XC4KVQ5
,[7]N[M]ZFC^RPZT4MObS?TZP/@Y/>2bc\GIeB&L6ZU5\:KQ]B(Dae7)<FPH@2>3
9@;H7>851=:a6KT+dG[W,:2P5f6Y:8YQZO&N35d8&K-BTeO:^8Ccc#Rg^L_f7;U)
Qe1/d9>CZS&0.+XAX8A5aB,1/5D:W>aOP(R0A[;S^4&5;#^SJ0gY:.Ja_)[<59&[
.H+[=W]4B#OSMZ3Y5XCfWaXR:QKG+aD/0>1UF\T;EX3gbH7U-CPT?W/b[?=4aN2>
(?(W/f>+RHHWHT;:0&K72/IUF_S8PW1De<fS;+AQD&5:6HG1DbMQ+9GU(F<X>&9b
)R0[VTX_cU2=V_7b4?-4EfR6DI\M<@.=KNSMFKJP#fC[/Y.f0Fe:(XNQ4db@aJKg
;3XXM3e@>L7FML;5]N]TRWMO&@4PAf+YHA:;&;/&cIVUK0E6SH^N;HUdWXK-:I/G
/Da6,BcGX9WPU5X2HJJ83Y9\H?#ZA]N@@f/]W6/+\PabG=V-eR5SDcBLWW#WD0#b
DecY-5/\;,&gV[M,LaS+S1[8CR,0AO8?HA,&>>HH=;QbM^_.D140+#Q35Z:F6NDF
VSL9TVFXF(gGW@69BJ=W&.-dD\cbVg,ZR.S:BMA-bJ1YCJ;0YPT;1OTBX4E#.K^+
:#+]9EQGEC\gfL)0/K^&DJb65IV+9COLZ5J,E6G<\RcFfH#c.2QVA(BFdP7I(/.1
^KLNS=AV5@U/\FQU=VRF7JJ>Y@9+/HU03U&;>W.G<#a(X-==^;f[YP;QO\eE-D7/
?DG;LF+_/_ANNYSXCf;MUL(cGPHYH[1HN?X&[1O5M^._<,0=.UHLA4JH7^X_88M+
XKf7g-0Q\];T=KQ>>F(02@/AfXP81I\VX]Q6]aT?e>WbLK6NRJTc^_BZ^DQ8=MAY
eQeWfX(<BVC0RVg+I7:0(+2Z=^9MQbdd7OLfO)F@CR3FT3&ZL9^I<a<WTa2If04R
7<f67S/FLM)B=I6[Y,I\1Y-S.45ZET=9+dIFH?B53A^\cH)XDG^,f9c#Ug8f>JFS
8J1QPLN++/[@.@(BE44V5;98T1@KNc[7&W5D-_]J;.NaZL3<<gb#PU3XD-gTaOJC
Z-R-eg=.=BI-;<78(^KFKMaUNT7e1(/2ae&FF@]RYEIUI-a[8=8:_TX-?L[V04GL
0g[-NF63R3,HZ0NeJB#8BUFM>:I>e1KY_8>WB4.GJ.MMPYUNaJ1bQKdc&35,FRdA
:99b7V@HJ^3GgUf9?P@>FON/bf5E4V.]/#.&/ZE-((4M<+/AE0WR/E_=/81H<#LP
McKX#Ke@gN.ZIH=3R?MV9K^gUG4:#)62[#YIL(eIaVda(/UWJ(>a8,GTVJEE[&be
,A_<dVCR9#5gHO]SX;A]\b:0.O70A_(V1S;YI.ZLDbJ4NDS2^7Ied/([=E0U?2(d
<_0>-@5CM(J\V?ETV[-F-2/_#9YQZ#6XQA@a,)<LbH3f=/gY6M;FFGN2>0JK2b[4
O(b>WT9^KO^9#9[ace?M@L2<b\ZS=42<5C:YM\21dLFR]IY/T?IXF\2=;5X@L)RG
4f[B-Q2>Y?];9ZG[FR0TT9MALTVU2EG\9b]>&Q#I7MKP]fc(_-#Sd1B_&R^=bZ6G
T[a5=FVB&-7E;OAQBH)4T0-\UXfRX8QI/eP1+DV:XcT@QFO4D7O82/XFO]bdQYgf
[N[^cKE4T:8AEaK+X?dO2>(S.6:cU8d9g(\TcZ_N+;/MF]XQ:F91/:JI0BC#BS1,
Q[Kc:A>_:a@TNKPS/bRb8GM=JFFRC(X_5US;BOLb;3X_ZZ);F<<,E+PO]A23]&[_
d\6U?=FMQAK@)F7/RJd(O6FQP<5bV#2EXTIF7\U]HH<CDc_#RL?71;g=\5H+SK^]
\?_-cMc&N>A:fa_Wc[UCfCL,B&Xg1HT\2(INDEKQ0J_KU)f-0+R7/&Y\f:ZEJ:AC
(G3daHK]DQbA87B9]PEYW#GWSV5#FC,&C:B?4DA+.E:Vf\Q1ebQdUeP/SAQ\YJf;
<bT;.Q3D:a9gJHf:&ab+LMW0U02EZ+R;RA-NXCP[2P6DRN+]1ZDU(BQNXHJSdH@a
Pf+GE@1e[/Pa5K#D>2GJ@a):D+TJ?be-N9M<K11fc#5FNQ:GZCEP.(7g:5X9McVT
d7V1/TR.RVNFEG5]=>#?^aD[]e,NTLBfZ^9)6<MBGYd;[W5a4^2+DI+#\DMS5D@Z
E^+;8X.01AP0PS.4dTA\,ceAf++C#\BbT[A[<bEDTN=@B^JZXE2YcNG@NV@&SSVQ
G7/E6GO&ScU/KK.Tb^W7RGJ9c]_PJBSBVC:8>]F8?VVGa.&[SX>VE]W/;5UGQ1ND
_T=DI<(#B.=0;:4g>43N0GSVV\X&NO/F;1+b-ZR)=H6\L,W8<Rbc+]:^]4:dV#N1
9.1\ENQ#c<.?^8#;9KcGE<U_7K]d\dZc;VDXgWE@Gbe-L;b2BI>CLc7J]HZa?cA?
C(BLV2:F);Lee80^[Y8^H_[4Z[8(1T8eOO4A0RDEg)#M5>b0W?SVf7IgccCTH0M,
P_H4A\WYKg.I4#(,B4\8L2.;Y+#J(Q.>fI^ZIQWO_824;+Y0^=0C6-d>e9/XW-?5
B<7E2@HeB5c5B1EIR93@(#<bYNHc+Q+RHK7(<&=ACJ=;<S@UBH/K]J2TB><^YYaS
7OL12MaRb0c>0PS4fd(g&)9<eDB^fUBN)B+fOL&(PUe_E>U.2g+Y3:/G&M<AAL8V
f\fEbXHEE)EJEM2V^D<D#QZ+/,&WHEG/A511c52Z=B&_XXCC\/6C/aNK2YA#K\6U
Y1.V-22[b,H+23K4E;W?);;]c.;]JJFZgZdX@HXGN8.UC_KSH+O[?UWL9[dUA@<;
3ND/)Y;99[4@E6fY^[._dVCb1TQ<D,_^Zc6GY;Q6/=fc20HGVaD9C=_aa)=3K0;b
W>EOY>A<98@9E2J/bZ,Jg-&FB\eF1F_3^6+g0TPF]E3_DeQ,(^CM55gF,Wf?#_UK
=_cG@TYYT4Md@H1FD,ZfTGN5d54]JX_>(24[T4]C3Y0:N.H\/79<SC1\AT]+e9RW
[K9X\=Z\7.D\[>M<ESZ-<4-C7cF83XGL5MT\fAV^6(-f)C/(?A&_209_?GK[RY#g
3&?71f3EU^.@?-:XR473I;[;K\#:Z07U.N+(3V&-,5J4N<Na,Q-4;c^KAP+bLfG(
2ER3Vc1N:&V(-Z+&UFUWV;35ZUL_738\(e6^JP]CLeZ#1[N[:eg>E4<,:LOX1(UG
.QJ@f5&.P-4=U=ASJTP;-T-/(TGG5HJWM19VYfaDCJSWS,?6b@=T9_1)=Me70@a[
=@Pff_<JZVAU8]d0<aCIP0gKP?5T1&]^[(U?UCH.5413Ua)R)2SS5;5,Dg\<A0P,
;aUYMaQ].,P]ZER30g?2VJ,;MLU,KK.LY-OIN)<IDNMf87OWK_10f;&a4\X_R;d4
)3TUdc53TeKaR/4f9P4N4-2EUgQJC.Z@#[K(_&R]F^\Pce]6P1#WZeY3Cb;aDP3R
gW9N.HbN@JU>HXV1^-BN>J3NbY+ABcG25ZY9PJ9JABPQVFg<\LK?2;V?\/,>,=^9
5_ECG3Ye>,H;J8K9=N&MI#=>=HSA81gC2#M2S/6XD0L#d>3/G9#8YK/Z:Jc(94W6
5.3&;Qc=5ZG74:EI(3,#+8He4?cC09Y7[)^?&=APO4[<D&/6)Kf0#A4Pcf:5&LD8
89528C?^4J(9()@EaGPd=B6<&I)_\C+3POBJ^_A,\e[g^7QC?D9ZJL2CT/805g)&
TPC#;eK=HOG@HM<E+E,6_,9>)+f(S7bF0<]dARXBTM5M))e:B1JLgV[bL]HHWE:6
cET0D(7UP66F<KG/C57TV4K5McUPQO<B8/CIB[7).,VU@d\@>=:eN;g]Dee^@GQ6
PPM,).K^K/?9?.<be->TPGM&&(c4G;cU#./YB7+R^d9LR[L7:^N;1[2-&(<B8AG_
[L,1ad1^f1(N:#P5DB+cV^NZ5LP[?IS>N1_geg]]Y:e[9S#dGA)&/0Dg:YaV^X?@
UX,9@/DL#:)=Nfb86R20/]9YE?NZ?Z:1BG8XS=T9>O(0]8&GC:7G6-W]6/;I0#/9
^Pc\),:.fbOFRDE=BNOfZKc@((+QCSX_a)GbJW?S@N1f8X@&:NBOZ[ODNA;]03=N
5(.44DJ4c8<D(&MJ:8FQ]_Q8AQ+@P;F?@42G9fD>0P/K>3V9fHQU)<1JQA-XG>CL
1,^5/#+FS9c2,LQ1V:O1b7:TRK,?/CAWXM0c^H;\f1-/KWC3W@:@bJXEY8IDRfSF
?.KdU7D(=JQGMaBOAGaKOb#C;C(Kfd747f?ZHYB&cKKeHITdYY-/LMIT6X&XV1T,
c#1f_&7Y5K4F76PS73,#ZR+43Fe/_ANFa656VYg9[@/dZJKUQK^=O4&ZI:LR.aQG
GZ5S437A)4^b#/^=48+EGM73_S0fVKWL7=X8HeK;^V/DX,48NB_(1bC\f^6#XbZ,
OD[?JBRE9TJ,MQ?(Z:8U5QEbS6c>/K?fN5HcP\TJCUKLD_A>7d1D)-,NE&YgVFTD
2A]K,g@H>dJS/8U4:LF-L:-2S(6a&MP5fHdJ9^^+Z>).8VOSOVCIW\;.&YWX1b<2
I_ZU2?g:N)3Y=XWXgEN8=e<bf8HW&B\+\F^EIB?)>[??CUa8GV214L6Ge5#X\_6=
&BN#5&D2U-(dPRV>/O8PPXNP6?7)6(0_BZ8_fN3PU;:X#HME8Yb;W;\^<KOa>Q(P
I;MR[08AL#Y-E^FeH:&C/VD3ET)4\(/H.R@HC8_T,ZReKCG&eYB1LI[9&=T+7AaE
Ia+K&cYK?P8R-2N:[JXH\f_>/,AMA,_@U?(^FXBH3:Tc^?P_:YXD7MGdSVI(eWWJ
)V1;?938<9CfRbWg5b76fI.HNM565EG.D()X2KM)49AcHCEM,HS5#&^(.Ue0E.=0
]5#Q+YAfNFXTYTNQ#]U+2&0=6VFE@0gC<:JP;C_^JaZK7#/&DFG\=#&=]c]J,La.
Y?:DM[e>Y2V>M4b>G\BB,B:BTKMEYE4Pa=U<Te@YSf?-ALE@:BA3c3L.C9W)28QQ
>DfCC[1e82\(4b+):OHRQ-a7e1]49@e@gYR?8RS@e[PJ6G?3]9-bYBJPWR+]MBI-
32[Q7=W__<04N,HIZ]:=1ZJ)8+a+2F_E;a@-2+5GJHeQCW_6WR#?71W3a96e<#\(
YSRVEL6eASH@.2C:H</6a^#-CG)-[N50_C=)V<RBM?J\^M/RY(fN++O_gFCOCS17
_+43:]EOc37V2-+]VK;b?_=[&(b5THXBd77LbaYY<L5c(<;8+IORJAe)_E;/Z(\W
.N&ed@g&_J:;XNPba6,7;6OE47O;::+Q^B)H?\^aSefITB<AF_=M]DK7M#U3J,A[
6OP<G;@daP-Z4-3OKcbT1I[Dcd_5b6IA4f=-5<f4TYNc>JV[P;8c,-\-;BEF-eQ&
:5>B=??U\)7c)_b]0[FO7C6:>HQ9M+>XC#e#C0>g\#T9LfZBJ?2c>#fAII31M]<3
EGR[;8@]C?KEDU?)Y-/BNYMTM9ge.=-N>I\K17OcbF;]QZ;Fa&K;QTUA5cdU_78#
Me\M8#(;\A+5Q3,CBQ6bg;PR;8R&1J?60ZDX3eHDAFHA=9C#a#)GcFPJB,_D_Ia9
6\SD0@V@M0F2:3@.X9O[gB(aG7\?daJ&Dd,,@_:=TR7&Z:c\SOM8e5A3JLLR@1-b
NBU1#)bC,?M1L\^Z&(Fb]@+WXC-USeWGNNJg;@a7e;c]2f&<Q/4]59bAbNg8@[#]
RN_\aJR>6A52-c6@T8.<9LIU)&I?c]Q^D6/Lc-_;LBgJGe-C&\:CW(D(->H5Pf\:
BW51V8V@,@[)a31:_.)FTUS@WJZ>[Od(KSN88ZOBgN4U[(O6e6&9@1;G@8c\?I9\
Q@/P#<6MYg8I/3LR<_R(1QDNc8,W4VF@A?)?XI)(c1Wce0/,ZNOF9dINKeaFaOOG
=9eX?cfU)(Sf1W6?M75HaHCK6UOQc0U^T]7J<4(U5bL1S:^?g]7^8M74/:=K<0B(
R0d[g]\>1(43123H?-NJ+.HM)C?P.2&+R#WV+>V0HaAbg37C-@27RJ4_ZF+KYf7Z
)]BU9@)GcAa(V,.FUJFCd-_[P45RDI0T;E<4\TALacJ]ad2@Z/-J7)U@f.C+(Z,_
PIaa3_0DVA2T;)dE,CEXPgCZ<OFXS95KLa-G438^GeB/-@ZL(5W=&LA7RJa@FaYP
K@,7.(K)F_4(MWNSX,L[DaQd:X+4X-7SW/bBaON>XV)-#3QI1f[=eT\@LF&S&d<C
WW;+9JKF]PH@eR5)4IW8&A2H-\E\8KFT4=(+>9C#U__-.Z2^,,CSO;S7V@IDEAf0
^#;37e=Ad2\_e[aIKfP_fGf\3TIe[_,YC?&[b8@F&CV?2Q[dCQ0.g/[\#3gXB]#V
4#3Z=YG@Z9V8c&gbBK.g8XDVRE(Z/a3KY=2L(2;bQ>HY\@@a>;5.f#)+d((99&Y_
OS=[gE6>3#C[PabG-,:QI.51,?MT0;OB=/0R?WYa&aP#=>G.6b#=/SGL24G<(6,9
cL,/1UMY.MSG+FcRe]D8RYBB:e>Te-,TA5g_HFSD<@WF6c#5:A=/F#814QX-#AX8
-9/OKS(YMd&KfAGM2\-M0)V)G62]WP14f^XYD9J5R0G2LXI=]58gZf4b8J0Z;L,e
-,64O2T-RURdG[-]fRLH<bf0RJJQ-^eZb0B@@P]g^bTL((/F[24&V][CcZ?,/VAd
8NK+I^XN<2:DNg-6,\N3XQe#\;]d3?SZ]BY8U&0DfA/<@2SD&:f]IJ+d,9/UDO^J
2gc/cGd^IFdd79=:/D2<_R>Af:3,J:W\S<F.H+Ve#RAXN<>710/R<@65);A2)/NH
>WOYae[5;cfEa.C><#G]&YUB=\(W9J_&<W1C\-4TI&FS=X-Y\10Ld/VWeT]>2<HD
).c93;I<@[9B)c_FLX0gTEW8^:Xa/8(/3[@\7O0532ER2)=fB)J-<0CF.Z[;)eTg
B;LFb.P54df]^S)@3EGOWJP:62I2[\JA]>MYQM/<M-gP0.5XCP#7_6;\f\[7XQ4)
;C/gCBYR5,IUa44Ng62X@W(MW39A7ZM/a&E)AZ=Y[,X2(5J6O)+f8+8ESP+<XF^V
gIg4-B@U9[gK?KM1^N?VG-J[+2Cb9+B;5N/<4VE#ZOF^cK1/F(],f04:N#T]KIIE
4bbO^3L&BWS?K4-<L.OBd<U\X\&/0PSM6DR,\1JcA(+B>;O58[<+](@WE)GG+RB&
V8e?>DYE6O^VJbXJ56Nb7)H6H>B/[aSO/,O?bNaa#XgQ0GcAQL\^9?:bGH3].P]M
5XBR2/SfO(8Jf:L\Z;3ESd5N2;S6#;F;e=K1@KKCb?22C>O.DTI]Ec0L4G\D@8,;
49b87(B26@fQ3S::R.A15(_d?-[D<R,Q@3@DAVC+ROgLB&MdB#R.1S((G6DJ^Lg0
Me12YC6&1fV<WaJ,<0a)Zad;)&^:8.;VR_,\TP=I]0T5RP3/FV@d\0_g2M?KAZP/
T(3>Wb\=[eED8Q>T)UH)0SJ.-?cR<+;Y:=O1_-/g3;R4[Xae)Vc]YTH7B-?&T)HG
KVM/A=Z[Be(>f,0\Z,L6]/6N.@A^Y7\7N7ROg\C-bQFN/&fd&<(5:BeN7UcF\F#D
G#<5ALLgV134RJ7J37XBeCgDZN=#+Ke_g>@+-#+_#-(L#6cZDX0PAJM4&]Vd4(Ea
3JYEed_#@H]NY4&94IGHJ6&G5I=;6/Ge,BQWTYVe&ST:EdMN]N9_.>gZg2&DK>YZ
;,TW-_0IW-D0dGcX7cI^7G4@4V0I55?eGT>S@X)cRK7XC(6IDJ\I,ZbIa8F5\,Z4
D3XPL5[?7:>POF-(,,XCJ<a0?2.B55)+1M?fe>T5YW#?#gb^9d^0E;EXTWVc^agD
EbQ]3HV7?LTC+7Q?6aJXT)RYRF#c6LPS-6#+[>)U=^#9J)Z)OT0(;K\bNIa<&6K8
)dB?=/86>5@@2(SR4VNAV(g9(X]bBJ>2TR]YWFM=]FR@1ZO=NRZ8\_8-PUS_G_#g
8R6cG(CO4(:J]#MfA72_E#Sg1Z-[E(B6GK-_\?Sa.OV;<6Z>A<QI0G7-+eL@-F;<
C#gV-ZZVVNG-HUS3L\AS+)&&Sb;e7ZU?/;eGT\(]2F?.#[17O51/>SNPTLc+5bS-
a64NdU#HYG(#)S8XF,-M78\4af^N=Y\@L<SKS9<?Id3;_f2P)QUTW)ES3R>):J;[
c;Q.VH.K&+3FPBV:KAM(<9>6IgBa/^^ADHHO+7ZCbZ=ZJ(GS?+AA7LP?a2M;fg.\
J_]2Y&;Id5-LL^?(-;@[V-T-7VH\N>,+4]G#AC/DP0FFab<AM=Z/B.Xe#\1XA\Z=
6e)RT5I#L4EM;+dAbLC7_H?[/S5BJ:3XA5UD?LTK0S+a>;,.;QS4X:cM?QIc.WJ;
#Bf68[BIG==e)+AdV5@R3/8cGd<ZZ([],b50b@8:ZJ&-+b<,.]:-d483O6N3(RYd
<,b-PR_T@W),(F&AZ0(-eQ50?4IgE^cHZM^^aV,QVe&SKV2.P2RMg1#R:-GU+5_#
^:C:B;I+\b+?gASa+SX/\6M?@(N8D2PDc51LZ/TTdQ@U62K>82ZPYO;Kf(.2@Q]-
;2T)5a6+PDf+VHZP\c3CRU5=M/SY:H(:,N5fN#0&\ec3OPS>9FX4JR.6<-TKeR,&
K8VW=:bTI#8aMa\PPBXADI6,1YTKTL^(56g/&HI>N;S6efH>&F.UcBfbQ.8H4A\B
><cGL0\YT-fA6f5&35(HT9OM&[J#1Q9L2;>=I3>\eT&>)f5J_MgX\OFFge[9Kc2)
3+Xd72S4J\ILASfGG=YRe[6=WUE7Ka>W(=/=^^,(IBH1(VQTG:ba/)U12<[-K.R_
#[3MZc<PM4c[g<R:Fe260[MIS;/&:F>JGa]UDLeC^M;=,0/E:+R<F+844OU;e>NB
\\g2+afGXC8Q7-/>T07^CgJN#BK+d=6-+0<-CBP<HPGd(BR8LXLYa/&8Oe>AC5UJ
?EOB([+,_(3HUPFZ_RVXAbU:8?cECd^gSINgIA#bM7f75BQ3Qc#N;b35,L8N10+0
gRH0=;FNESCG/6IbSKBb&Oa8(#56dD+gX=LD2QcZV0Y1e#,gKZW_8]:E@&NeBX#?
B,NEC5@A+;\Ag\Z]Z/LR/I-+,NMSD9Q4DH]cI^E7G7&WdC0ZWY=D7843CI\;6WT/
XgER6T6b[[;L)7P.K_.9NH3._d9:WG+&2<>S?#-G7^O9)P)Sc1;T0))2&dUVXg^e
8VFB^9PZC0_QIAI#1)WBD]FKF,Zf\9eWM5<5ADHJJ<L1ULCFNG.]I#4R#Yac)(EC
P:Z]-RFRdJ7Nf\O=@WFC[eYP7I7^A/+WPeDaC;aAUYS_bT:<VI4(&=<6:GCc7,;^
\=67R_@g.Z(01&<M?g9NWLZ8SB)>=2&Zg89-gJKgB[)X8-Y_D<XbNYS=8RQ0:Rf/
8La[O)0QP@:)U(;-.LJR-_B<Y.&OI9/A2JWK<MQ):F8WVV2.)?\,WSF5I,K89HGc
MJ#Y3ZPOJD(aYDG:g;U(,=XZ.B[>ZG6c4])K2Z#6gH0[NUJ@c#4?&K<8(FB-ZLQB
1g)=cR#ZH^36eY74d^F8+G9BEUJSG&_MbaB;0.4I>AAbE>ga\]MO^7fLBU3f[6Rb
)#]IYZQ-E3Q4?fEM:]NT,&84>Q6D3Q<D6(6?<fg^2LBT)\,B=B[?\/TO\^.>EW4,
\fe:H>U&0KCe]bE<>Cf[G^@)]<Ha0;7e3f<Q]f9Y,>bBW4?B7eRLfCPb(Ff1_fD8
c.TbXSTffI2;0d31[SZWg6USQd<TL(X]PT8+f#:b]2Hae>(Q<Hg;,6=HEc9&+RI\
DQf?gY?JT2IX?>YP>:UO4W\WY\(7)W#\>ZJ^7\>N9b5X&2[d.@V1E_,JAcS#A79H
[+WTPSW;::Q<Ha\0G6J4\fDg<WFYY739VbG+54ea0E#RdBC[.<GPT1b43W.TZ1,g
=]#aY-#B&eX,M_dGSX?EUMf69e?U[365:+>3S(@IW.8Vdb<H.I0\<79c1Q-.#QR5
fa6,[S\K4E]LFg_.Ob^[)T.fYg=F@CPPF#XAD+dF+:4SBOQ16,];/AdBaJWIe&&A
&a6,&aRcA+2D+O3:930T6]ZG(ZKOIXY?1B@087=BHK:WXTKAfNaZQ7>Yea,gNK4A
Ac8\<U4.LH3#V/6Wc&O=eH+Mbc4-PCYE1.UX(-.-/D</HZX?=\C7Y9V-BKb0>8;7
>FX\;V<I&85.A3#cC5QNNR3fU5@Q]B&_=Hd.9F;DEf\+DIU045]DTNJ.U-2_-7=P
I#;JF_VYN&ULdg+\I3?O6V,=>3EWD,0KXA+)(D^;=9_/6O&E4(6RgF/5C?H:D#:\
R>=]<O37Oe0gYc4_;]G/\ORW^=>A4<-2RUPF,M@4>07\7GML0U\Q/<16XefX=ZUT
QIR8(9OZM8[IMHQ\Q#7?,2d(EbZ?\/CCY?MU_]&5=J6[-Z-(2Q[Zg72P(DG1X10>
[58,_5J05Y,TEAfX<=42(6F5PaRZV[-]R[bC6=,PD=Ya+>(3N#f]W[(;\@VFW,2<
Y2-,e,K/2KVB<]P3XMBG>X-D,WIH6>5Q?F,I92M,4XULJ[//?1J^39D8\Y^C(faA
E>b4IFJ751:#0bVN94e0/SW7c4;02LKOBRFH\A=OCY_1]:7Q1#/MQL^IOD@c0/N^
M^P?S5<UMQHU3?M5N/Bf8[/\13\Q.Z0JJVG\eQ_&@JFPTW9@gfHOMd@C12DRE[#Y
Y4PRB=:V]dNB_2D65B0<KJ5fE;_7XW=5-J@#g&W;B+Q8UA:e2H\PgKJ86K_<0WTX
M<>X+2N8Z2dZD:AOFV+NO/)_S>O9R1^^JFYJ<G^Tdf^]YDL:dY0ZPSD#:5@T[cCQ
I\Hc=,2+fcDKUIdF^<:5R\1bb@,&G7SEXQ77HU&cfVeA)^)^g;Y2SL^M)6+<5gd[
\BG8N#/RCM+CX,@dN-I)A^Ie-,C^8=K(AG,J#YE(G&()V_YK+6WLYO]g,OJ3N<M,
18efD_MESWUTeNJ6VNV8@?V(.N(P>DXe/_05E\3dGW(f84BM9GWWL,,WYXI(c(g/
T\>eOIB8B@XAcLJ4_<?B397@\Q;&<F,0,.?2:A&]=RD#MPc.<Pe#PL/R(^aR=.ND
8WY964,VOORY_7F,PJe6<#,cHf1=_NYYGW4T?A]e?\Kd2W#2ZE3)[3G4V[K5FX>8
1Jf4=HJM:=Cg1I)ad;)#bAgg3M:-FQ0E99G<_V?\390Gf)>aIe0,J^3[G(_#>T;V
H754b.(06\gP-G,>GYQbD-b8KM[/^FQ_KFXT^T#aOO33b\;&LXOQgN9<^.IZ)]a.
,dV63,b^=2I)=Kd-]V>[LW-fb()(H7@W)bR3T2fSb0)Vf3L]B>D,eQD.LbJf57\5
N>881MB4H[=Sg&FU,TK)IB698d.,[0F;ZI68\<5M^W9aC/<68UHg+X]F,A;R72@Y
PA]Tg;H>&Q[Z\717D8/4EET)_XT\=>I+W&PNQ^YN<)S5c959Z-7dA7==L:)YF:CX
+A+I9@]7aY2O[g;a)<N#6D_T]</2U[c#FUR_>.E(E_2T6YN9b&JgN1WE_3E57^eH
<b[\ZK.&F&MAF&^/CN7R-.+047,0:C\g@XPKTa2SSVWJ0+&[ZY>TC5K20H(0WUfA
XN7+@LZEd++c5dAF38d4VR;;XZ]507NA+>\]<\G0-LaCe05\6+aZ_7^PX.bR2-8P
P<E^,>[5)KH(G.O]8]4J?gYG0+Hf;G#d?b@B163C,-f;Vec3A^A0B>IdUPM<HLJ(
5]:KDcR-9Hb^]-.gI9<d8:B[5]Y.b/aGMMKF]EP>YaT-1KY/C04KW/QAFFIZHgTW
+F5,A55eQE8WS_>_.9bdTN5S^9FL2JgY3dCg::8LFeK]W3--Tf>(7WACaeP#D)[I
N<W>+&@=BM1)AVfM[LG)aP6<,.)X7,3>-)7[#>PLg;ZeYJdXL@A18A&_JSQPB+GQ
Y)II,/=R9agT]\XUTY,_N470_M9FYWM]BP)D/=&DAD\1_Y3.J2b\fbdd\I7_9Y_/
7+9RcG<.Y6G<+c:XM^XTQWC>U-,f&PU/_==?e1(-RNO#76>N0/T;e)bP[S<U>S<3
E)DZL#]P>bCaWQ-A=,3W/IPNPRC8P#@76]75f)^6H59,DKJF:.Q4-dZTMZEL-f4N
^477R6Y^-TP46]/0I:0gNSb\JZ:6GQ/,JR<C92^;_HZ/N>3/ZO843;X#[ZL=/GF(
P#.HDLR_2VE0UM=W(?=^+T-DE:0VgI#Z[OYW.E]IdWGP7[Af.^[I_PB,MQ80bR#Q
P<M>RC#dI8X]]&:6B>f/W<cA+HOO-Le[56V&[APdV38FAH9g45ge5GI8KQT[&OPd
+c]N5+0Y]ObMBbOeJVYH]b/#T@eL8Yag\K]Y/#_RU,G5#V25,->Mgb=&;3Vd501O
c&Db2Ued=;>_b-O3ROagPcJ/Z:4HH)e,:)/>[,-beK_g4R<WfcaEJSb@-5..S#J3
GN>Jcd=T.6)#e7/d6L+?_.#:[ccFK:f(Z->\UT8aRg&4e/G.A?SKVS4b:2c:INCF
J[7H[J4d8AERDgKYT>NE:P88,KIHV1-e)ITU2J(KI^Lc@V_:UcUEPDJ9O=68J83U
F,f+YgTDAO;/,ZUEY=Z1A=BbJ112-7FLR/YC6<c<cV-1HT6GPccCF[_aV]cJ+D:&
d)-IM.Y/7Kf^NY4(RGV#b...AQdIf=E:cA)]b_eXRI^911C&GI>^2/I8FVeWO_S&
T)@DBM2?NK01_ZcO@1)I1CfAYQN\^1[PbbG>a)/HbSBQQ7MD-V@\0^ED2S20YZ2T
I32RW8ObDI+;G=,S@A_&]=9-O(6,;\[4B3)^b6NE_]XN<FO>7[@6(8dMUe^,TB(0
aI5J;[CX:?E,c0(e6/V.6=7gSS1_R[Y9UADSM<?ZF@0dIH)\.E1W3Z3,)1/^YNXC
XIB1A;;MI?1P1G6f-1WGb#:A^^gN/S3;ZLVN0IS<(^@.6::N87F;3GGH#21fgCcN
)/7^WeHD@0RWHX0:_:#P<N1Me-#/EJ]A;Kb9:O].Z]ROEW:\XM5:6Qb&,ZD9N=OY
/S.U6QMEUf@gLQ6S(bI+MF.:Z_[UP?A<GT1;_>7UC+bW\VBQ/W+&6Jc#AfSAf.Q?
]<Y=7J;8&7TL=1SAEAQX#;U-:V:U[?LF+KUB?NggE0L&--0-&M;)=^)5SCdYO6,M
4.UUJ1@B-D=g@1fN:4cF4cf-7:-2+M.EcB+J.LebSU;1H5\4DGCSBP.#g\/bdFKT
H(?6WB?XTYOag3YLeZQc9-9YR@B,VW4\#&YE6A366W^]M@CJVZ59>>7]TIJ/A+FT
QB]Mg/@d18>9=XGU@24P->;WPMW2AZSgK8e)W;bHB;U:N?VR\=AJ#=V4<FIU#E(f
O@.AD_A;c<R6eCB&b;U6=dQ_M?&>BB<^e,9>)Jc0BOa(E<FXG0XGgQKHg1L)-44U
)F]DKPDG<@[b@_f6eB6&F#-;d)a.OZMa38-I,UfS4OCf[R#;ZR++fOe1Q4NVC>0Y
eSdQd>D\3(2CH0\2BZADHcX-fT0cNAFg_0CHT<]4[7D:])OaC(^?@N1,^L\5cC9>
CHR:+13(MSJ>BV&(^TaN0.^-4E(F18&_DV6>S,58KTR\Y]O]8H5E@K^+dR1-^G(P
U6ZL6345BHg_#=.2&]H1(K&bW+4CaPO\W)YW=c#aJ3LYJRP72UOT5SNL4(KeX+fM
0TM6?GQH]MQ7cI)SZ@5#,>Y0BBLNb6aQ(/Y]A\?<&<WU#?Hg-OZAGFU7RO[9[\9A
WY]0c><]E=1g-7U9M/V:&TZ75c/_;E#Ca8/?)O,6(HVeY3=/C^/87^a(JOG(X15.
EY5GR-[M>M35O.H@a,H(W6Z_8S,RZ.#]g>,8c1V-CPNL=O9>Vb,B=N@3Q:3-)c)K
5YW;Cb-ZaBaCgLe#^,PaQ92db_52P#f&=-,[4-f_\6M9>@^d,M4Y[.AU3+Xe]6G<
#84+OM[@3TcZ)T<4[M?]e7&7ga9)^RbA.XL(.O_O#MYc],d_(cGEDR</)Q(-IQZ+
G#G;UeXS/(Oe>GH]FfTR\LMd+E58Ec-I\eX=0a0^G.QgaRR-Oe@Z@Z?Z_cCVU^8+
(Y?HD9]dGC+;G.6IDR\JO7R9GSf,eR6[YK&G0g3QOf(.Jb21_]fVcJ&:37]+0UNc
);]S:IDB@Y0g16a19)c/2;eL;cJOFYeT99S_+(c-#K-8J\?YA#c68-c9@X(2Fd_=
HTJUIBM0SN?M7ePTZ:0#fO3:4.6YE4E9?eR;.LF_8CWcG[0-VF0=470C>O5,><A4
.=9E>[&+:P,gNcMZaT8NF=+4XAU?2EDc6J:+7_.YVa3894LD<#HEYU3SSY:@gO)1
?7S1;Z-)T)<K[b39);K<JN=FY;Kd7M4WI:P:<9CUI8b?SQ.<GGGe+3L<+&5I:]UR
d=MOFQ8G.)9.P/O:/JCPg]41-.9a-#gOY9\)_^/T8Q[VO[U3R@#U=_O.,Q.R.^)W
g/(^H5AF(1/dBZ,,0JY(DG@583]=/D;)V\5&7W9=9,/G3=R@>;F>LXFN&2)XV5QZ
^?7:ZE4e?Hf5MIA0;,Jb=cYA;_a6g5,NVTF0HT=)Q\^]\//91cHf/3#JB.TGMBfL
+V#^S8(Z2IPd+VPfXPgHadM03V,2Q_<1M)?KY)dY](1:YRNV-7RIWPbM_4GL#[WW
.0#NX]6#9a6LeaA:3f[WRd]FJ5^K-0(JF@&FF3FX3,?GS2Dd,9#NPH2#&70SP=+e
/SZgW@[2X19gcGWU+/X<JG4Y42/,NAdQP+f<@bIgY^5T34.ECg@&9Ie[G^#_OR5^
Y2RgU0>4/34]He6.b@I3g=\\.7cM-6#NZ;9,4K^GUDO-f2cECQS/=?#R-=KX]c(9
8aHLeD(4/1?c+5M=1^F.Lg2/<FR4E6?a)<<T[7H9IJd;gCgA4OEcG00-[b4#P:]_
1Zf[;:.e??3?1WV.SS8?HA6[#0bNK-cGMXK<2S0RRHR\8<R7R)T^@G?dL9&=^aDO
-.S(gB&,PWFHL?@Dg4)ZaLNaDF^FVf(H2::,.gV)?>5GA\6WY_dZ/1d4fVeH]/U2
,OeA[1EUD8KK;Q=?D<(88-)HW(HJg-5/,^FHX,+ASZG:U>]cT<\fab=#XUea=4DI
2&.5VdbR6DP.=4+aWa0?:]]L,F;>d(aIe=Fe^0,M7PK+<WW(0>F=>bJf+G/ZB\ZA
H#B8(bVW6QXY:__CHYcJP#OLW5Mb/;TaOR8d2X8(MGLU0=)49MU;?bJ8QHWU0bUO
2^TD/18(JA)Y)$
`endprotected
endmodule