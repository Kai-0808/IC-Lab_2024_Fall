//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
oPCHwnZfwvpVBvv/eyC59S29oKsOZU/V2C1IJKDHXAf3ZHsV/4rkD/GvBFFt+Nz0
MbcNBelgG8D/+jNYHFd3FnwOoDJ3+KC3zqGlfcJiRvu1XhBX2cOPAcMCT8c6QsJ7
5nIWfisrNj40ystg+62+pz/2xen2USYVAuZrkW9tUaPyZv/NJdPG5AkuiQnfuOuA
dq4ARdL9WROLRAG8HvDFmZmfIU5wG4zbM/Lo69lUp4398PCQN3rcgHkOEcPx3wqP
vSqsKgZQF6Svs3Qy7OqDv9g0LSxh16Oi7TAnD/+YakornVYsanhVtABr3rTJBSGe
wsIYHXoVFXB2O88iyTPhMg==
//pragma protect end_key_block
//pragma protect digest_block
o7Qubf5bKSGYrBIM1C5xD/T5pvg=
//pragma protect end_digest_block
//pragma protect data_block
0R3oDnTSlMvWBDJB8JhLiz8atsK3RZFnPDWJ0KA0MpnJ+TD6OWAp0NGHr/zXHxTO
nN02w6asTbcZIWM8aTFF3+HQx4JCoSfioht/1/5AyzrjrcH/BLUfYkGeudFOdgra
ahLyU3x2Tnonx65MZamKRvKDlilEhBrlYj9sicahFejWkSN1cu5yvCIF6lxYib8I
UWjH6+E8pP//9yIuZQ1pj0rqlh3reDlmvhXlQzNMu4nzx+XT3SjRs/Q3oEy1RwqL
UUf2xWpijT/YEDeNv9s6mYs6Stau6kZogB9BqqmO6p4ljLkiRAimyc584LBLwf5n
qrzVmqf5tCUJJicyBsFNiF9iNNyEJjTgJdmCPKAQUN5QtxfnANLKfg3XQSMZIwCB
mPIrIuqp27tXzL5ujUyxnf/93z0Cjnr7k+58yfgURctXfnPQcyNoiARJlPW7jt0/
2uMSlxX2iEmv+XPt447xHg==
//pragma protect end_data_block
//pragma protect digest_block
ezsDXoqpfYi5RZOh6l0YCNtZInY=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype.sv"
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
S+kn709brJba8cKulV/fVX8uFov/PXubIiG/zYBQuJJc1lvbV8dkgTqBLWv6NBJp
9Mj5iwEbidSsvKCNvba08GhKnyCovqMpmiKHCkmTqP+6P56JQEuFbPMQBpL+kGDC
w2VrvsQFOn/p/TKH4oAp25AK9+JCb/zyQDlorGsUMI2gBTgI3Pp6ZD7R81zbiO6W
TVt+ybZjVZo5vlW03bGVvqBMKFy7IDli6mVg2a920GeLIG+C/ofwXWEte3gbh2UK
zRIeZ5CIhDuS2Zomj7d0DVcd8cOgqe1tzLJ6E7CfaoE1CPrY+XWsmsjZK/8DqGp4
DSpl86sDFUZ0poEimX6H6g==
//pragma protect end_key_block
//pragma protect digest_block
4jkWf32T+Zr0cBI8t3K8p9lH+x4=
//pragma protect end_digest_block
//pragma protect data_block
nmBg4jIh1UcpKAfSWmj2C4f5IH5rjjC2aTzVxK7MmeSj6G4zhalQgYcAG5qH1iDA
6YQ0s/aN02NZIFEW9UAVwpQ2rNMbiH4pWsKLR9LVAVP450A+qSSe3q9pqdtaTnU5
gndpbcNaBFIV/Updfc2iOzuat2jixPmWszQsU7JDMmK4a05+8rgF5kkyGAnng7w2
uXumPcPZVxaBRHiNzmvlFYlJWP2YBXSZXzlnfSVenfwx/KATjIoIn15O0XgPGoDi
dXJ+C2mka9IvXNYTmlwBYubC/gq6OsW4vdHLpFrSHmHLHH8E/duFU1ZftQQSv2qK
B5h8ZQmEz8XaUuaBmgvNxro3GDyjw411TOZTNB9kT+j6cDeyEuknZtATwc8/Jara
Zcc+7d0+zkujPj3XBbAk447Kuj0X7MBN378P0a07zMCDyhhM1ibj8zRuXicC0OnQ
FFzqtYx+Yy+Lwzc26LwtORqf+WSxKGYhhwr+SIcB80EDr/6FsP2VPB6nPvuuQOAg
8zomXhOftfBr9rIidjzDQGYdf4weEY7V2iucPFF71OjcQKcfXrCNvM8uMvULmjUF
o9aXFAcFYeop5qX1ldrmalL2txF4EroPxScK3lypNrMbg8H26iUsMdU1ItBgnuSN
b1/T1+c9VlBPwevK5ceVSqPTYTzjEasSJrWHOFs14VppfTbf28BT/1Zk86DONDrE
kMq4N28qCxTa92doUv5GFYPdmh18z8FsqZNg2pTg9dfsZ6tUB932mI/UOKvtFuKM
M4mX3vjnCs3W5dPAs4FaBCYtIa+UYXDOOJr16n61OInZcJlTmQWny7ahee4tHidt
UmihrYYNRahlODhI1tM5gVjoCJuBnKCtCKMDm5yashFSH121pmFIYKKGr3b64FSY
Z9fXvSrtqXGnW5T2WVGPJW4HbocOZzB7vTfcVK8UZ9ibiuT9M1l4VUh/5QeRQ2op
1Nogs1TX8c+fJycw8kCEAtD5WkwxD7RC6BkCbWyAHDLP34GOo/fuVvsCmepSu9GB
PzN48dyWdNsdMFXe4tjOqsf3qjc0kqgZbZXutbxqWTL2TJocrLYiiPIOm7nvo0lh
T7InONx9Y2HMiPRVtBnh/KBYFxcttd7Rl1Hrr08kMiKRKl8BHgrI3dBW0TNOO/a3
AoATPwSmGkgivpXULdYcZnbCjb3oF9vQ+1qN2txFVtMmjyKV99iqCcaozN+TMk7U
3UURMAOBvsr2noeHFcK7zd8xOT7e0xr8P85OdXwR2wWT8JFRzmLe8KKL5Wga7KgH
m1mJguq1/A3ENUqSrRsGuLEQ+9/l6MjbfavyFQ9GNZIXS+qqKvVRglreWNxrlGh9
d+9yr9JL4D1iEiHrQom6H4qrNUbPehV2HKeIRhEmF0rrXySTE73kevJm103m9pYI
trRahK5RfRAlBJUyG/zV3QXO/H06M8LfjRLTkYnUNeL5XOzqjq1aZytvn5GyqxSb
52yl0H1QE/m41tZPhGRWA4Uma/PB9HqFKXpTNVoVdnA/gbY5XEkCXDmf7c+EGhsy
643caF2vkoywGnjvFotr7c3uyXw5ag9P/sJancJyLKs7WBH5rWJt4w7Bsd/9uZ3+
V3H73nGhE71Ej0TL4Fe7NYaYO6tsTLkUCq4kyF6ZS6yJCubaDBJnn461PUBkoEvi
TMM671lqcSpgFzbhv5dlAM1BUsQXTX5NprX5083pFXZ80Z2O0m7jeGZJqrJ5AV6x
EHpHm//pgNxUiqtu4v2JEhrPY+NJvF0XBNVaZrRAGop0AJwIvPF7fEMbVvjcif6A
BRACow5paADll/qlbDu0+zQEugulCJsuYSdnA9o5k5TsV54uRW7bHsZxEydsFGpm
mK8VO1WQ5ZS+n4LxhwXCj3tcmDcQeLnRV7sx7n7YA6D1oRTp1Tr6nlIMrshkzqf7
DszFvBOb/j6CbaqWAFB/PZuhduPV0U0c34p5axKsgmckoW/X0qajZ2IgXPweA7pm
4E/KiR/8Xi/E9LtGUFb2KgxBInRHfQu4CZzgL/UrkAJM0ukX0MVIOxnA3gZWAX2o
+IPX6c2yfangdWKm++RwvLAJJ0eyzGi00UnFY341yMYt0dD6rfaw86txQwdFgUco
pVVJ3r8Pz7FmEiA2NHbBC6aidW6gbKNtS07uKSqsirodh8JMTnf5Q9V2GmrxnaPo
kGEw5Qk/G2h0RpSbhOAbeAVScyX/i0kquWvv8Jev+l2cRI7PN1jgrYeKDM8JqXyr
yMusMjlSAq9U5nghkN2r4Hpk57442PNUoJdc5Y8Jln7KvelogpB1C2uXFl16Bd3d
KK5kyQ2qQpzLBDx2SIrFziL00RNjsyuR2M8qqwmrgIoEThEL2dnaYOdIdmte2rOV
t+7EvJULiV5bbtUEI68ZPDMLTjVdEwYZ6uAPRweMU+Es37gltvIgwaTcnRBb8Br8
Vj4GhQMXmKd6553ruBDawlfvEQ7T2LyHwD2oEKMjpNNBUpzHytdOvNtSSLW9ckg6
AI74PeIrfdVXaaPw+kqIsvICJCUNSV4tXfWV9y1f8omCukjQwYVdSOUzAXnkaIm7
rAAmLZF2MNDPiCQZ6bFmVtk+aCTFtaaN5Lia3IqwW0uZ1/ec+H1ERB0FPm9bHfMp
59PFYlGIp7IMFIqlZ6/lKaWZ7Xd8+kVtukgzWSIRHPIjcfN1JmnI/kiLWEUoa33x
PPYtmYWeNEGoZ2wMNB6VGAdqbBfrz+FqSn55Wvmyo4oSU0gLEpDkKpWNbNvjLtKR
QckQw0SmWVBuNXjUR9VyFA30zpOaIZJ5hNs2vkn5b9k6N4CAZf1tgWPZUfZikmun
ThjwGPCdWTO/nnGIIT3F7wrOO+7GPwRFdo1YZd3r4SRPDyJPWzvlEGxgsMaYo/xm
qFmvVlf87ssFYSzo/aY4S0ieVaithVpsQY+yjczex7OPp0sYsDNstl92A5bA/RbD
GZckjVtcTV9poLTwYlxoNbPIImn+JzF4BKWtS6YgffTpVOCeySuX5p0tGra6ZNB7
rxcvhQC1gcK44SexFbtbTbteWVWiOf3ZRq+44fQGb3t8PAyFcq2crrtO4qXasXkY
q+WS+MezGUGIk5TZseCgSr8fFeWhLpgIJ5F3ADHokrit+nfKAM4eJQB7j2Zd21O+
KxCi5BKMQvJbHp6jHyM/Vtrlm03FPzinPxM4J5KaRomTPEgl4XiCpgU57NH1Oyc9
zWfakkNHFeRlek8EZS0lRrPLhQRM4KF49J3yJLApIzu1xgYYdAsP3XQZDVKWkWuT
pUETDCzf+CSTn0jeiuEqDGDAuwPzpDpx5N/46C2TM+tj7Ulmfkzgqnr6DsheNYEW
S4yVo4dTqHZemUhlsPX2xmDC+Q9rl+Zs/gwsg3N8ndvKWAF4QTHHurArwRc2jdjA
dOxqXHObiu5cSLOEgdd2GP7hIshtVCOKihYrD11jq3D0ENFDixUWOBOOlQFIxN63
tBDCOdhKXoWF80if5Bxs3VCM90ekI2+b+hh3OndOsumK24pUxUySZ3k7eHj9npWU
ZW1djfzlslf/mfp9OpoW5u7gg/n33+z3nopdSKJQr2liX9xbSzhCyQptbWH5mqi5
ePHclB5L7yl55cfO/UC61Sy0fnaeIynplTU7ckQZ5ujHUc3aCUXdYJw5bMKRt4rK
yxMUv7F5oa4B7yuL/EYu8UGlXueeq/WpldrIAULCwTuzjJvUe4UjhySILwYFqMfS
J38Ikr4S83v+mWsWjP9z1tbHkgTxUZCQtqzuRHz4B4pMHHers6AXV6b7oVUqBf9E
61debFkFsPshpdbhhP75TBMkPEFScmovrj6FPiyqzfH53aqAqcv70HmUHf/X8OLz
rn1wNee3jKZh6eHBOca/lxhJChQVwL1TmiXIq/MsdRoxkOvxFw4KuwILHMj25DRw
zsGP7z7oZhRQcg87UP7LaWLlodStyC70OY+AXJxjxGpyzrzso6ms/kryXz4yTcxm
7qVaoRno43LtdScVwc+gz4fCS7AjxuL2P87e9BNcmBt+Lt3PTL1BsxWrDxgvBr9A
2ICM0A0QfIkzYgJgjwnOp9WM0xv8vTpa+u/OuLp06A9J1vbL0uerHmm2msqIghti
sy3zPBCfwj9HwqWxi1HEZuFcvXGQsXqXek3sg2Z9DYsicK8OzjqmqjyXFivOfaN2
rhIkxdajTGvivozriABoxPI/DDIar9tl/84qRDsV7FshZAKjSbuyA6cWo7IuWOgx
U9yIw7NaFhjqZk3Zy8KIsNaQY2PKU0ly6u/dXwtZadX97On1UAABi83HKDIV6I7p
HlGQit6E28ja/TxnE38g5ktrnG7p9gpYFFJ4pLZCrjdoTlag4N8FcJTLGKWK26RY
BmnvXG3O3aiScTZB+d+YRCub+KwIIKoKCe3uKQnWo1VbqYupqJC8qs94e//XZHP/
nX5JFNblSZL1UK+nV4dL/DzazWI3EigKdtzts+mMCB8ivHmj9+aDvWK1KNXV2jic
+w15WJNZBL9ARKFVjnyiViV2uhsz5vBCVXzckrHpQJW6LGzRUYzo/89fNUNBoItd
jTTPqEQV4xv5phY1VtDxyqh80NFkuLrlWYcsnBoNYoV2osoyMEmcTwPRYC1ikfQa
Ygq2VKwjtpzyfrpd6/3zrE7heezmO+HwGTgNTl4jAAY+uPuBJT+GCTfwFNbdMdP5
gF8PPxYIMOr2biDaXHvp/skhFChljpY2qCchmNAyl4POklV0iXXYDimAYOhftVFo
JnYDhts/3WSd6Rc/Mt7ljI+XCZ1kflCo2BojQIRdKSQcFcqGIbGrOYO6fYLfQMhk
loHVEkpj+CPDaK8cOvloQQY2nWDK4XmPLZGoPaspoyaHV1v67+YrqnT7/lYCg56Z
4aE24ZpPDLLlpEXPZoDD7kD0Gb9NvtB9s8LgrInHysn7L2Mjq0VsDjarr1Wltn3s
BKFSQSew/KGGqO7PdN/2OxsqDgPTyu3eWUbb+F8FPEKtKt6OnmbHMj1iEYcZIVNn
h4FZzGQikkpuSkL991nWtAQKEtUL4Bl0DOHWPOvk/sFzxYiiYYS9meQa5yVjqTcg
Qzo5gwIRw/Yh9AZPPkH6HQCtMom32axpjMEPyqO7h7LAAM2LoKr9WLMg0Kdu5/P/
z3SsPtc1MDLohktGSzzpx3MnwmsSSSVULIoJY85CI6A7KY22flMiQwosUaB3klzq
y4l35XeYFFitLAHLEsDr9j/g5EQrnUB9ziDjwlFautRJApHcURgTMJc4ItoBeDBQ
ZngHXQyw8opjkDXOK/95BY3hhei6+f7QqRrK75rDTjVVhl2k+WwKWOqiGazFD/wf
34et0e/g+kE9FZR94iDg26/YSZKtwPUAmfpzwMbfxaIN5qPFmp/WB1V42vDzE0PS
0PP3uRe8wAe37IaKe1x0h17R14BYMHt8PhBI4n5cmPiMNb1rcmG9v7tVrl7QhNh/
e6o80L+d1Ir7X/HKtL+W2z9REiJ+NWZJlLQY/M3P2qD9Eni3szhLFQ8zr56XPzD3
shv3T44oZoclPShaEqH7y6tqGkAbioJWPHI0qfpP6uT/HEiLaYmQvhSORkKIaF7r
2Ls7gGXs1h9ofqHJzLj7M4eJ7Mh0WJglpfnIicfco+VHws9hhU1pENyTIiLlSx94
xHhjI/G7Iel3iWcnTv0GPR5/hiskHKhWErXdmkdg5rT7/b/dmnidQi7ak8Lfdo9i
c8WgnyNkpCITb8zg29ziwsP5LZiAx/no5QPmqO/MGHAzO3srft4FqyHuuGxwFj5X
cK4/DcG7mRv0ZEK+jVfdJjSV5wNHlpu62JzB956kjVv9KYvoMmxVkMMCDYjeDvDT
rsu0XQwUEmoraBfzvt4x9QKaPk9WdrcCljIwGt0KqhZiimeIXdiYzKfKH92XQgU0
PBZwiAT/yyhvnVC+FTnTkWnrt+/hOLDwcQQFgzKQZM132h0RRC3q1Nfadw46Rhph
DfXH8l3qzfIi2rOfjKy9UXKploHe1G6spGLDp+sEv0NzBEoyd4Y1OkMJZGmn1Ncb
DaXdSW3chGcyr0F2ywTkB+L81rxEcBtizLJsSIOvN8CMLT3Jx4ClHupVI5aP0Ji6
l7dLLhTIeqwr7RM1A9OngNJ5fYy8pLP1DihC11dKU/MSlSSVQ6HRhfqiz5zxawnf
FJyxINxLJ7dTpngHuBaMqC2fo3hGVV9DrcbxxDpU+0yEOGqZwNlovT8YpmjyvyTq
sWt/enk6Umc5v9Wv+SqUl1F9nSTBOjuXlnE4tgNP91daAoxQ5oQ3RNpzwei7GwWS
iIY2/8BJfypUBkewdnWF8ENwz+M4gNGeput5+j3Lr6k/fKXmenBLNhAa4551SQSz
dUAV4gFG/wpBGMhZ+WAuN5oO9XcEVz+kcjoJ1emIji/gZ2yXMpyXzWsgFlD5jK1P
dpRdXb5L8spDI1sydP4srQ83Cb+sBabww7qGI5UZJjsKxgKXhKp0eaW3d5rMUKLN
lCndZCz51S/wT6WFzNhb3nG5XdF+0J2jTAT/IR1XOD+m7tc7paHyLlzvptkfr1+G
5AJrQqPkB5f3TWoR8duRfrV+1ghyw4gl3ZO3qo9fX8gownXmKUIPfvm9qJVQyGA8
9bp3riHCyhmFRHxy70CryTiP7hfkhZgey5LfK03jraM6GW5zvgyGuIWPK8JLJNSf
Y7OBrH85qjOrmgG9JILSKIwqObd+050YcPEORmIdw1s1bw6pTxVhPMwHiHA5MkuU
jhYX/OqsGwAs7dvozCWPZhGKmcsSyzrRXBSSZnlmFaInb6pIIZ4+AVBcvxUsXMMI
dAvadsCyVNpplrCI38VDB7OjsBULyK3YKAEURaXqqUD9uR0ehoI2Tdf5MHjPdDJv
+NX2zQJ+nZPQ8d9cCG8avWmzXPg5Zgfu5cWOBYUQCpOzNVJBwXGnS0WH/T27vMak
f507Olxj5Bj5TFxvo+XISnT6xpa/iFK3ilaqEFTjocmLC4Noaw3iJd8ilKK4FBES
01qMEwUB0yIqUH+gmzDF/eqL0Lv1Huu5fIhKII9CRU8fOt1juhs18EqMVUk08QR3
zABEHJQCuByukmOgkQqLR3zadGm80OmwQmsgZQ7R1E+dKGuHBKRnVZy3Geow6ilW
dq5URCC9rsz/m4prWejW61bfqZTVH3wlyaPnFt7ACIOfe4YMab1Zk9c94S0ibsJ8
1IhwlyjPeDcQyDLcFo7GWj/AU7sfdoSbMnDk5hbRyxmiFd6tWQQmbMeBNNTTeu8m
v3OfPocvyEiLu+T20myhN9DIY94FEh8UoCDXJSiA3JrJkVReeSI3dyTsS70rEXAo
FnaXH7zYrU0ops40MsWrupaDBM6LUCo3295rVDGER6Y6NjcKAxmsqidB5lnYixhQ
3Tr5vjm+3g+Dt/blu6jDKKN5tkRtyCevh6Zj2W+45DKmJX0/ywYJezR6VsT0E3ni
Qta0B2ZQK093fEZW/VL73ZBtLaq58bH9HklX74dX39klFkPN/QnBSgKL6G60b75I
i1fMcNLExbtyVepGwapJS+ImF+SX/4p8bk+vcN3exj4svYyXq6aa16EKBChP2owX
JhL7BH1NQqSYM4tptDtVB96Llf6pjxu+c/1ZJRLbNANMqnQwG8DdhZTYPLPlUz8w
e/UKwJmD1JEvhOvfmJLzEmIFO0SkJHhYvwSx5mekh38oTrCe7dRoNU7x10syzD0f
5GnnOoz+ZywK6zu2gb8rZ5Qulw4pnqv1y3uxOYCFBvhvMyxIXjPvOfZh6G91Rdy2
Nz/KX0WIi2MIrFFju/5MsqiT3zDwGGG8EoLSk3ARIcnXfUUDqPRK3+Gi1CtLJahH
yWd2noZd1MDjOx3C6gs/5UhNmK7UtIUejieZtfpXcryT0QZQRK079tw2yxLFYElC
Ym9ma1iXciLOQ6TxMQ7yTPqVjhvx+g3naWDM0OKkVyGXb42ItJ6aUf6qfMrU4wPL
vT8b8wgIo8GqB337eMPz39sNrdNCJKaEr/AYrW20Roebxsdaetc3oxf/SeUwCjVP
2w/eY4Z9PmSpWetS0oMJ61zmPYxbhUGm1alw6Svqm3/LsHbGLLBJ9wKw4Gsqr3xA
VCiapQN+uTKfTAxyjkmmyjciMvIKt2dTiO/cqApvuPImm7qI328ED/0Xh8IZdhgQ
u9iWzne59znRtWXILPZwlMbMTOXSOw3IpEyDWRiO7pKnWTliePhL+EYvaVibW8kw
lXRn/51uikgfzKal7zo4cgovL8AbDYDMRYyXinTkvP0DYPDk4b1k+9i4+N+vxDyR
i5/ev6AwJIMrPZGxWxl6iL9IWOc8oDedWDMHUVUTjkQzFIajdX7Z4r0tTzU1zR9Z
0tO4UYgeFbtPGXRgXLhs5emBL1gqG3O8nlh1vSWrih8N7g/5/OMZi50+n8JqVC3O
OvPPQaPdiqD1PV0nYY1BUW2NWbU8kwl32/2H5ChpMLRjiZyofS5o49mOd73rtEAq
Lg3NgpM9oak9dzpuW0gweNQ2YTgYd1zmueQBNMXxFNeJPa44Pci88Yu/FluiTtBF
M0rXxwVs7qV7vIRqBkodsCtVpRJCY5iS994I/JZPRJ7kSGUMADUb/x5xuiQIe+Bk
AhmsGzyjgJ8wZwuEPg28adt6Zfg097XjuRDwtYF/+023TTF57Z2R9FR2NGpGRMxv
qWMssmcbO06Io3EHcK0qWSYNZzUFStpnDZQKpIAaO8BEVV/DPN9apHlALS1aPw6S
JbAar6XUB7ZlqbDs6dp3OpoJkBHWycZqZ8O357Ett4wL9DUdWbltwmj4+U1PbteR
mvMgf3RtuBkaRdheBPmZ3IFH25lu0WivcUl+Yitcg+m5RvAl5fOwBiDlTwHCrpxI
CAZg9zgPTtqdRM+EsQ88bHSMb5OnDlPOnzcwKYDGa607R0ZPhfB9s3AAMHuG42g0
x4AMYuZitATDrdy1RdLb3Me17LnxJKOtl4bn1iSLTMyW+AdGmxQXNwlliVbjYsul
ye/addbvDc7QGfuyQP5jd/xkCs06LsFWsAJReefmDIBC95vfxkjyHrdGZhD5JiZr
OeiTpVygiJa3M/kLKTZNGUrL23NNsYpN1vK8NCp497U+R/tOInLg+c/N04HWRn/i
sr0V9+MaOWevd4nyy/T9nqFlHt7jI0Zt7o3NGUOnquG3p8i9FyfhWRkBMDhIWo1L
/laW7LXeVyksNiNSsLNgEBW35H7LSdw6fZc63r+N5AXatV6xV6tHHaomG7431lXe
0H/dtfi/nrVEvVZ+bYnv+8jhoTcRZ2JLlt8/K0nA+b7YP5b46NSAgq6AzukX6qjV
LNyPKNEHdbbQFTo8CInU7hyz6XJmDcw+npZ2Lxk1kviO1TW+DxZVvp/ZbpNZL1Fd
kl1ZQy9wRI632TEAEkG5yDZeH/71JQcTB/sO9YvsqajpedoFZTnDeIz7ekxRWvC+
iHZYLAgtRCwvtDJtkv8Y1QKC1Ng4s7BzoTuk5eqniSL8CDkFMnHNRRQm1tQWO5UI
o5uo9NsgiVZzhPO1c6Qp7J9J+56/+8R0SrNl+OOURJE5VgLYP3VuR7in7lfT/nXa
coYRZS1sDtH8PUAV3/6f43CIGFMAvEhgKziyu6Q41CneiHEPcUd3Af/S2BtDNu+p
k7iqv2+GJVKdvV/AFJ32i5Y5r92vt26hCKWcXljDMkAxzMkdXhd8qlrfAPwEXLmh
78saG67uJkp4/4+1jn4pK1xgdOywj4RT9vvrSTtIC8gdta4ELCvj0iQ20Vp8W8WU
Y83M22t92gyVClotvM1e9GyqVNfnQ/ks3VXMUQJh//y/dLNnmggF7ivHazUfF5w7
vqeLxQtsP8Yaj0CIqoadezFeJ9+79oUf0Egoq2Fq0GaDmURa36eB5J7568vKToKI
nk/bNhJtLvFYKwfCd+hpzVs4eb4nO0/VYiyRNakEuJPK+7f7Rm3MIMmjs0Ul7Tjl
bdZ42RK4xVS029VfyPclm8LV9xqklq1Fj2Uk+6wsPPgWe1Teus/BGIrbP0vCV8UP
5AGxDjbmBjG14C9W+qwYGP7++7EeveigyHcEhJhJS3cz8K+5ztwW38c+xd1afqkn
F+rhOfJuXxejRGwqTLDLE3uFxTztpeja+y0vk0ViobgZfkNf/9C65/68+R+2TZR6
t4rLrZPmH7R/OxCLzoaQ7Px3MHYwGnw7P6wNLfn2jVtaqb5H+F/aOvqRn8EUTRGm
+FpVThzixKi3JjeKrtvaDAWQ/aG7oCKSthYDcJ7tA+TJ8lKJE0HsH6B7N2PYYHI5
0idXpV9FjVgTICDkdaITtrR94DZ8JI68c2c/8tlSO+xMYUwtN0cn26Rv6o0gj7vC
4R4vW2sXz8m311wRjyTy+pGMN/RzzAVkuOrkem7+G6ysL+mBWtj+ZkSL4SejFw6d
erHVaFjzOj7Xa5avQFUuNzZWelVp8a8Kkm2cv2BsgM9zdaUFITprLSGqwIk1KaNc
Hv7A6ALbTMp1EawZ5EAbDSYIT3ldx29mImWvthXQT63JF116eQ1op7Oz0lk2I0HS
kTdcOXErRMpSZKYv783cOUVij4OexyuPElFgLnH8JCNlgntvxrdEGK+EFsp7K6Mh
31bvp33uUHYCwwmuPIuDJ5shzfXAHi0yElp4/s+c/Jp0JgqvRSbgzlcLuT6LjqMq
hAvd5JUN/dsL1KModRhxMBReiTRZ3N1/1tfjEbCIKQB/RY2KuHsQkZnna6kyRB9A
PhXSHMXnA65iS73m2nbPezxOZC1dl2N5JpCT5pDEW+HCmcwP/+wysWGWveYLZpjY
Syi4X8zt00zVB9+kzqlueEfbRdt/RvE6Rfk6WOVK1IrAjrx0MO+us4LGyoPzzkpa
oP/V5ne9G4RcrBwcuizE26rFBgHvWXVdSdweaKqGB2HKJXb7zd00FikjcONzOOjV
paJx2yCR9MPhjeAey8lUwqhVbSduQZuir9xb0RzzDkb5ZuON0su+KloLYzMwX2Xt
ahMScME6G69y3hr2+U4TpdFksDGRCik8QJTk4d1ptVn0wna3lhbZBU15iAfkPvLC
HAHWAp06s4es90WiS3x2dbekAovDorzxsFbXqxxtg6roFSqdsTnI+zzNDQhwwpRP
UPfKFpJmUfO3a3Xi0356+9cmjLcGvofd1pguQS9CFkGldMf3fqC4YkMZLhM2k3rO
yrO6LkD/ESG1TUfOrGKHCBaHxLSY3txUOUz21g55lAw94TtFKkSbstXo2VTUa6Wx
BWSWarKE4MHB+XNP86kPeEaV4U08NGTRxEAfKcaJOH4/qrN4/JRdu87UU3WgqAyI
5YgUC++gq0l5ViHtrh9eu1LngvDZi0zudf1lqI5jvtHErfMxhGUHmq0QWG5TkUfT
EBBwm6lsj+txcf1oA7M9sAG4oiTo5BCvIvhXA/omeiz1BnHcpiwTuELV1eVhB2JC
AI6LF+D0nDrPnnUU/Yu1SWT6m+aq7v6O1i4mLr0RElP0fz7kUWd3WqEYvG8Yj6FK
YliHZioiQZMWb5sytwuUgiHwQn0OxHqQCq6u8Cy6IbWf/f0yyu4wf1ypwTBuvU4h
V5qlHAJle06qxMxo/EfC8CRLce3tEG3unka/rNixW6pGE7jT6+L9u5q9gmtMkpxo
fx/YQLiJUzybadxuxyWK5VVD9hCdLhTIWxtjBfhkMvMor/aXhB3QGFYaFxLcbiLF
wJdIryW4yLJ3CQInT7PCa2BzIACA6uaofHBNeVIZ44dn/cCnu2SdejMfChxkTMSm
UdtMbPOg2l9jJXj7PzqoLfFqWgD/Hqk1Umo2Is5wGlQaFY1ZUBhq+OfahjCWpYFZ
L2oxtNYJhiTLdNiUY/VLt32f0XUbatDpbTmlVTORu+JgA8T+9jJWv04EqZdec7a/
J+VDwOb0knsep+/W1lYRQXsjFDQc7rWXqQWPDE0F8PQtm4OxxDTek5+ZcIJUUpfl
FyA7nOnJoEaizP15eLLco1ihvXTBhoRXfyEA17jt54vJO4I9Dr8Mc44vj+HxNEEz
MMYlYVNr2QL0d2T0ukCg5hCEwyBE0ILQ5QMQLo8lKA8D2hA0fNUdnDwptaqq6n2S
YcipnelqJVO7csEfNQRDougD96zkrgsZZ/jSFMAZsXFPZrBjoqQECOeb8TcozfhP
L70ktb23e1sRzIdngGaMAQQ8VE6gcgb2jQkj6AhQbrIGVBrFSTOwHmt0F/LsRJ6a
fsnjrhEYaehUK6pwnsdE02AuU+mBoSn+6L6wcF2Mjdm0/I9eyEVlXxCCjDJKW96v
ElpPq0l11J73g8yh4aT5q7peID+ac45M3fTgYp7QMDPykY5ybaiXR6hY2BQR87MY
GGhj4Bktxojq0lmlQcafvAdoNOYRLWOn2BFNaEG+gnlKGUgexAWSf8IVffcwbAcg
BiRFMGeAYDePzps7kg+QWC+wGo8IHazJMXU1RDic1SgLVDrAJT12YgIRxoT1fKB3
OtVQFcWm0PVV0HIxxJ1IEh1nllhs7eljv8vLQD0KQNLWGEy//HN0Ut1atE/SK5+e
vOD2SAmiPDqAfD0/VwFpUcp5kk3dWQ+Y339YhPHSF+YYYM3LBenaEKSBAVlzdAvT
QSXVF4OQlEmNrk24IPKNSjx5IMmJVrDaLBu/YmZoMM1GrPr0hKfISebqm9bNz6WY
7Je32OcXF/UHrkD9LXBdk/GzYq5k8+pwY4gLot18b2769x72HwjznRE0+Z+j/CFW
hTuXUj0mCR+AJylJjyLkcMNc9D5cZx1kZXyCvhBtdhaZtws4NnZf46rKm7m0EyLW
3kCl+eEVIyHEmRhxi2gOIHefjYHw2K4kQr4VRl38hk0ZnUpef4e+7Xi8HGwWN7FU
ROtON4xXliKF7ii9lXbWgoR94xru0K3ddJXRan8KLui4OPOEUadeQTUSn8ISoPes
Tdmbo+SsCWkIfgR3FoZLSM4tOLqckQfxvcjwaG9yCEXrQarJg8hzyzNK5u5+qcMO
ZFMPC2qC1XnSQpeq3k9GtLoparlKRbylWUfXcqCzxxWBsZp5Ll6mrpsWyYPSfbPG
OhNaGFpCVFHHF5Yo5iVlEfkWHabeMAzdd30PYdeFSjphq9VmDgVwIA2QqeWNk1Rp
vhIhjk30ARU/nknClVFpp6WcgkfzQ4WF5GdB2FXPWuC1GD/BAQd+ERoe3uHTx2SH
50r6x5JCPp/qZHknY0P6lyoV7aPOSOXxEO9IVi9OCmKGn4o4oBw+e3CiKAbf7g9J
F19ry1T+Y4QY7fGXb4+WSLOqp1lHsIkrpS1iWJCH6gBvMt0aN+A/q/SOq+hLOVYF
EacP3lg+FwhaALOaYO1jFxN/DGvfMINO5cxLixg3suRoEeEMeIUVyS6jREbRbVso
UPbBSXjfKztsX777FlvipqwaBfB3JJocei8cOXlsUGr0a3xsX0frVnZBd5LgHkkd
74pMREw+YfWpGOxfgeEAd2XotJg/CC74aC6h7DYyOM+HsuBblmwGIo60tDaZsFWp
hNs4oBcQ2v7Rs8sgkUbZTdpMMFmhvs2lh7X/loY2wWLgJEkXaef9imU5nm4xMIZ+
RCkcGv3piclZHVmfe+cyYdsF2ggrNYvtc8mNbvtO1Y63MmOsSWry+/8EQfSBCaos
CP0QTSNcHpAiuqhDNBLxtI4FBvyoLRff4sTEbDy1XuPjQTpTfjlnXNHFPv1Aq+y0
2Debn3uuBl6A5TzIpWMF9g7JWfZ5na2iu7keGxIlweLIBTTXmiLEqRKqpJy/H084
ahNMNECMd9q2PrtEPpzCo3f9EJVgf7fOw4NkX1PKE4Gh8NLosQcqvh8Uxwkly7pG
SOyAOJMWG/7Ne5rO74Rs5q8yIeWuMGe16St337m7K2lRRw2S/N5FGanx9R45Cl/z
8+AulRQpkP3TwlOIyXWxaG810bOK1oLC9hK3S9z+x6j3ArLzX2y8zTCvRmU9JsKb
naCiNhAy0TzqME2dtj475H68nhfWEc/62zuWQUygpj2ovvyAhnAVpdD96r70RdIt
mEgc0e2v1QZZ0fG5rdhQ7+K5R/LreUfCl6oQ8J9XKJLhFJS4KJSiSgStLOGa+GZs
vjNtSYDxfmLQ3Tf/9QExaLjpBlJGex+siLgSepyeV1M6W8eRIw90xaedvaNgXnyB
/sj2gyxczeMGaM7LsYMvkJ1xG+XogHgjvlQRRm1ol1iQPtB7aqeTLYUdK916oMk8
Vo/ZREIZ0y5MS0eXkpDE1tqA3uQNvf1vR9Az/IkYPVxqh6IU0g2ZEmTf8eTHTVcW
fHhQiLIozhygdmZCa0w3vcCmo4vuXOZJcyOxd1R34h7GiWjYVQeS5DSwnyz7NeY/
fq912Wnn6hhcc07eMlk1jC92JeNPHJ/cogy+JDB9XWhXSe0uWDoP/6HvkjJT5/9s
nOFkA9+yMyBsKSTcm/tdtMED/26274nYQVhQGtpp7Mku4Vh/CKN76t8/W4ALf4iI
LSHeSTBAV08FbAZkCDmPzxvngtKntsz101o5F5jQuP3fjcim6g3Ok1xj6CHkcnWe
dinm4F+zZdP7RErVhSD56bkCtX0lCRm1HkbXBpd4INt4SK+kZ0AmUnr7aIWIaona
f7TTXoPw76ddZAdhyqXtmpbivrGffh7OUpfuIDINQiASqFayml0rlH8P9RX6u/7L
hBfAL+wr5U33Al4I29djXOWEs5F5oBz1vE3wx7SsAAHVu/Tu9DOKK5gxvKCCynCl
dJktddt90RV93EwZG4o1oExJsBHbzck27kkLpVptutFR+zJlabRQHFLb+OVth3W4
5xS7H8sgF70gpuVjzv1Z8cZ2EOksjcTaCIYvZrwRVJR1tCYohSZgJa1l1ZWL4uJK
jLIjtKvB8yqDiHaBC9IkV5KgQm4bD0FFSuzmV1zNbE4vC1OBDyUNtW2MJYflX1cR
YosXddr5UaegFIvUC3oP598imT3hGr6xY3KnJAkDTtUPLUTc8tmj+MRQCIoEr1Lt
lfCRAPTF3s69nynSOqo5aWyNcgzhbPwSvu/rdu44ZlQzY89dZuXAltsT3BWrf0l3
ep8uJIqLV1usZAmyKTd+gnM1brFEnbWqre+KRAmS/9Qgq7TRTvUzBaHK+GETjDnm
tVDb+wsGlgSO7aoAc667v2MzdZQtwGyekdPMN7ihLB+BrVrYfotK3Fm4QyIhDZ6v
v7uOf+XswMF7B1A+G428K5PEwiQQU8Ql8/LCgaFRRp6D9YeQ83A6n6rgXLCn+ZxQ
aaBF1/w2n17PTN30w2bY2B4PCAzAYuA80FaiQXp6bryvNr+5K4fkkm/wghE+mzpT
0H12mVABUhf4/RV5iUvM8P/NnT1FXjcX/JJsTqji8t31ONwlpXOi7QSSkx4Pwx5v
pitzuiDuqxoNYcQsEevZephABqzLMBxiM6B2ad3XCmWrUxDFdK684AefoivGUT+7
xAQaSfQZS4MSiVjJ98itabfzcfNa6Z/AQKZ2WeTSp5+1iIKzZOLWIa2fjmwa/K95
xIh7+W0aor+BtMqHjt9znyEK0E1UzJBjN4RaQ1ygDj16u0JvVuMDyWC3Pfg3Z/nV
rQPeQOYErXx6BBvJNM0yChNNzMVtdRIn1LafzuysYa+TxzlN/gZ+tKWO3YElJUms
dCuLAI7NMkxnawupu8sIizAlfSPdP/LVB4sRboRrR/zrX4+w6LomFvf5/L43YnMD
QswCNc2TouFsdHcN8+z7MXgirEIGXRyXSkli7+FmZVac4OaFErnZw2gYQ9Q/eBMg
kZ5tfd8i9eLHj/66BDRH4TjY9pbU0kk7uIFw4lJAwHv2q0rc4zh2PgGWc96hPDKk
AmMILsYUUBHKiC0uVesYwQBJ60NyREhvUKK5wKWqg3jSNTAOuGxNdUz4CGq4jHmG
ZHuKjJS3O4+I8+sig8w0gqhSzsV0TY6fiejSvkLzX7/9BZEG6Pe+UBoPew0kCbPl
Zd+raWwage1RHJf9XOAYunQ4+MeoPR5SFbrf1DS45AgGJ7NKSwlUH9+GLmwDIrHu
QYMD5ckAujJg6ISZL5I+ddQwnVDU55MYLA9DqjldWsme0KQ8kD+Z4pup49hMvLFK
QvaICeqtFxfxho/FLw7A68yNBoLENj/UwcQBqiektMrq4oV8CfbzqvIxSVauaZ6m
ZIVlB8euyRPWb2pdt7hht6izguTkFGR+i5+qp+nhX6IWD+vluoIdZNghSsGujlmM
+79hvgBOSvr5oGawYNAYNoHVT4CwcpTrQ+33O53BWo9w40GzOXYlp6Mo6tF7iEOv
n/r7CmrqSmOk7A7Tn9xF1S/r+t52zn1xTtvFSVKkv5I3ih/u31ubKVak1KvqH9YP
ViV+oQfiL/BRnT8xFRlKnzFycxPWZIeDoZZGXe/yM/6XG9zOUg9Oiqvk3K7945yA
BgH7Gt/k0v4PQgc0g506w4mC4xjPQOjTgNZ0gTXY0RCN+YqB3fK0FYMFgvjrk4nr
DzTDG+WIGvpoCE95882CLcNTei3CE1norx2Hifh5o2fijKOOG/uhWSs62zR+q4H4
ZKj/mXTjPEYl1auNNugPxai+upyyX71xjbFArGdRV8YMcqEiI1lkYC4QwyOYPqYj
Eyw0NOdn52GSjt/wj1PJ40FfKgNJ1uFcL2ssV/MnsYOSCUB27eRsPAiqc4BfWwYt
bcwgEtilLBtScvbhIDHE5zMlcxCleM6AW80jt9aiu9WflOqJZiu7UPZMd3uy7FYf
YZge9ONb2XV52tr4ul9PuAjlwok0kD2sOuL5y+cd6/z23hO7HjHsYeIgSlEtITHj
4UhHollVb0KNVyaU9cKkH4i9NxVbcf6Qucuk66xQmMFa9CzIIlWThfbVvJ6ZVN8e
pOonsPzSgrJ5zRNcl58bVUO772NjmQQTo2CQfEr7uzAS5akiTM2MUnoyaxwIecp1
KOkKDCGaRdeobsNO/fVnV5qAtCspTj4czxvvGzarMAZwEqNzrQnqtPuG9DmQdlMV
41FDtnNZMZBMfgCa+Q5VwnSZiWXVc/fPaC4oGl4sbxpjxexBIp3963g+nToXlMPj
7K7b608LGXl4Swb1XvRGooNmx9ajSlsr03+yHr6p0AdStUZSOvwQx+s4fO7LYjsC
Z5eE7IS1URVbejS0hYbOfZual+hDr/v1g/1I70ZpXYSLt3vp5+xJeT+SBgqiGsdP
Y/fIP2Qlr92BjT5ag5oultadPX0Qgnm5agNDql6H+SHwoLhNZPMtHnIQf5dlDm7U
j+vKx7NqoiHpPsvi3CRhGnu1g0uZoMKhA6z5YvIFI8dp3CHBohpC+RB025djmOkD
1FoBEjieU/V4TqeOpyQvNOQGMtHKNt9fg4loDYSodzjGVAqESHhWuxjgMoJy+GQ6
26kmHy4JCnvKUl4k+NrFuk7hslW7XYowxlajVngkJzdR3wNkmo9/9groLWRoYUWD
RF8Ia59JHFUY4z4nyFIHO2A7SJAyF5/3NyIJtN+7u79SOCJdwd4anhlmOGphdqM8
UQLZYP0/MugJIwkDsh9UZ8iGzhPj5asFhIOMag/YOOCuWzFnBiUZWb8u3570Aw3A
QD6OxCHXYYoBrDA3NFrmfFvLTGzlSmKwtMzmb+q6sU6AfSDjSxrv7LHENzSapsZt
cOgOgFK6ISYKC8HTruTYcpz+nZXYEau4N9ZEH9VNTLXHC7joFrMC4WAlHAiCs2Or
VygFYfK0+/mVR+dr6ZGjopRiZoZxXLylAk5VQkKWgoPmrRwMXpFZNLf+aHPN/x0n
hBraMdUYMElyZ+1rPL9JaGkGhQCLIhfyqkwnko5kBXNFzwXwN/rVBL1zylA9JOjq
1Z6FDqSsFfe99rQvLHmXRPFkTkC+zG8KKm0X+BJ3UrOfyMB6KaW6NylkblatKbr4
ezmeTsi8cMBT1QrHPBLovvIKwGR91NGlXZompGREcwwLp/5BJ2h/Lsnh4abAjZ+Z
ffqpLki86OVvoQJ/zIURonOVsoMyr00gIm83p3S66i9sRNi50L/O0jAwgUDuMFbD
r1//faSAhQlq7tlnjd0pex3aM5TSqDhgufBPhf3Olhiugk7sP+5K1z1T8ZGFAecw
X+doXWwKG3vlm40WYE1xE0VfOCOVexXeR+4/g39KsBOaLSBMhJWxX18mzG7uv4Vz
RfG03dwHRVhtsr20t9MwnjMByffA8Hvc2WNuOJo8FzwlB6276avj9Uy5KxntAXfx
K54gRYTxCPpaIW8ntvLmaqKYlLcEgj5QKnnoV7RfWxM1BY40LsaIecmfHEWYs5dc
L+ZSPVGb/IRM6zYtlHiuaqJzO3RXSA/i0N13PUEQC0ueHBbKBFdK73RAsGDF+RqN
NO/WQsMAP6HwKBTtrmru+eu3obBSkoAwHrjvSs1M4oWov6aI4keRxs+NCLzbh9s2
u0MfqWCQsrgsVyQiqbumd24GycvZ5/f/G+C4EXeEKCmCmXfKUGtqdkDM3sppbNJw
rDUxf8WEWlTlPaSzav3iquMxzjxApsWNYcOUQ2fdV5Un24QssV4f2sZKM/QLnB5T
pOL6uKkMEq4qJTBCqpyBg684rI9vlNowb31b5JQLXTuwYElMd3N2+PZu69uqAM+O
cOapw/6evL6aPARWKinU1iboxN1ebH4o7hRfwKMEk4GScrw6YzRWFwnEoMdOiPS7
xAEEs9TAUR4Gl13rsaJZnDjkZFhIEvZ0Hti1ug3EuwMfiRhqFS6etdudxZAGYpG3
CRHWdHzCZuii8UVLTA3oQZ5JxqF/4+v5ohGVeQ/8uLod///jGUIhUw+V/s2oMLJY
CGAXPD9065Np45KTE3eyLndLBEsC00GVTtpFq+VW0lHAOLytk9fShZdFFVEfqgHn
Jg0lsBWuGkaBuqV8/VaSmyTGjrVOecOQ4cGMWOEO6nUfOKQaa3y1Vj4eyOQ1T8qS
NEMCqt0s51CLmWmyPbyMI1X3atxyhaaOjTSiDUXpVh2GQijOxWFdOco34hxawYZi
jTySYXGgS5CoEALvwgHYCtK2Sch5vaDQk0JCNyw3Bv5q7Bg2iMcM8kV8b0LelfMT
tYLV/2QFXlfck9DQgBBi68dEk0/YjDHlhVu6wG8BFwlLFF1yH4UoGGCcCKuP5cBZ
AsaWvk+MrqyBWIqHZ7gSsR4qcPhwXu4c8D2RjZH5Xg7MauUtKr8H3QBSTWjVMTOs
sCH/2BctSe3WJZIP3406IeA56Hmxyp+LHcOZMgv4azZ5KVU3Vm9W/7MO6Pbhlnbq
ZAgVl9wN2GWZpjk/VENrWs2jjnpAxf++am4uBiAOdSGMp6ffyqKE6caYJW1e8ftX
EfamL54EV44uRWffbOQwzl0e7jaAehid6PNQB8PR9+RuJBH5WDqRytbqH6gItkYB
n5+B7/KvqMhSQ6yd3LMRB075H+d0TNrRO9wbtLVoRVmZJAje4q7kGeLn/FEDID9P
nkz5yIa/Bszn/nlsAdZtIKgnxo5x8BpstboHSrS03TjZ3ih5/jJLBWyUXuA2Wcp/
fR4tesj5j/P3at360duMvp4rXG/kF7Tvxgdx5z6cJXZL6NwOCrkMI/HXmKfPccbc
gO8Vi4PRfxTD4vkDCvWt4I8Ta/6v+yHHvLUKMRCbp0itWia3xJ/qF+gdPylYY4MB
eEb0s9k/D7jo39ewXtZYSDcBkdPUy51QTgMCgcRWeepN7FLmrgp2h0F01vKwZySw
DG/83KrFri6oSrZFPkXdwxUTJTd9e0KlIt4emoBHkBAnKePNS/jY3eTAw/6eiOpf
9CnpZLgzuLdrQ0iebP/xq3lybf0kTv9s6WM32OTsn5xoWZUHad1wzWGi58cqM7dh
go41OIvS/0LEF4K6vPVfmNdDvWWTJSXMdwj7Kw00eUrC+m8M7Ix/QcovCuW8hvte
wv/UDFLOHZAYmW7XrV+Nz+jKCIs8GajyvPEz2y0C5t9Xip1uZxIl4tuDOOQtKAuN
cR3TNfaixcFf43BekcZYlFenBXBV+q2KXXhm8t863MKC12H4j5qlrVSYS86rrg+J
Ko8DWZgfFc0QPV6Je57+0p7u7X/V9UohNypz33A1RnoJiCDcBognNztAicwKm/16
nrg9P33G0d9TGknD8aHzijRyaBQ9i5Y1QvIG670ZwHT8qJvzYXIznS1yWTjOqdwn
YSz8hllJfNzGBZn/ldIcSjxGI7FxNr6RgAEjbQ0ctHz2mYjqrfrfldVm//pJNDp7
XgILK62arQyBJ2904I4PTF9u5xIybI6Fw72Udu7WSH5xOhzBramokVirxKHjinz+
ZS6ml+j1v+u+QVbXh4rkSg8xUECgZIKbzo5yEdqaoT9mhFfdfQpNhPBs03iyQqV+
eySePy/V6uVjA6tRAc5LBCsGREqjwu5+L2bn9mCanc/ICJZaUhHN9iSBAF1lWBaT
kiU5TZmWyubjJFm12fsQu8TSIgmgc7GSQiJ8h4Yoo/eGg5zVXTa/F3mLRlTkZW4/
bPCDLL5s65w/vlNOKoR7yCe8upGCHORP/bIc6OacEq3danPdawokM96WA8Ft69FL
fbq8TJiY5ultT0/+57c6fPNk333niNTmkuvJ3vdnBVuLLwiX1MDEAotsDh3OtZKf
BAYyw1ZpmhvCuFYQIMfREF0+7I/O9tRDd9DPHmO78R+0FQc+MJcr0V/mQ9dJnhSb
Iu6z6e8fA4sJva+otWME/osV2V/YdRJxpJDdUeisxmuYdBaD0WE/7KxiNVGICS1V
1Px6UGxlLEhJCX+HAtbkf5Arti7k7mRQ1q111CuN8DP7ZU+9nsagkPzw0ublDGQt
sc84UNTnUkN+k6s911WL+C0zzZy43rI1TZaHojauj6CZztzCK4qojGOa+s0lKXL/
bFMI5vLEphYkxkxjgttkXjNYA03cFfn7Itr0UAXuUtSfXD9Rc2RzHRCaVHkvKGbm
RFJgmpmZmFcY5+8hdpIydiWUb3Z7m2ThxZC+uVSdNhyPdd8WkP2XZjoAEn5VkqkN
2KhbPmL9vfqDRVynklrjcVQY5jf7nEZM+FGwOjAeEaboN4SJnJDYwzEQckiWalEE
KZFUvF/kWYJh7DjUxN0+cVfeka8WNbZ0EPFuCpYJfiNe4s2T22fS6g9ICbbZqyTm
eLvtVU2xxJnTIDNzGYP+R5buHcxTP6fOX4ner9STYlEaXlYNnW2BBiu5uAzxihfr
IIeZAGGpneo2tsuCpbe/akrFfBZ6BRMAspfkNKn3wgpX5B7QOCtNSbPfTUH85Yua
C7nhIiguko9zQtaSBMpwk0SGj9SuDX7Jhqgx9SHtaOUWOkuSPQoGAHkmRKER+6h2
myRKKMEb9/8MWHxOlhL5hLtuP5GqNHwWRoxTnV7+0zxxDZ/gGMUPyKd1PfLPq5Vc
9V6hdO8IyP5MDlEwNFrNZJxWrAYy9bD/TgR47RUsZfgbFLSC6OOLIDT2lzvhQVFZ
VWbAOx/8JN5neTvXR822N1cGuDkcx5w0Nn+TaSt2Tks85eGSWy385gHa2de68gtc
x7CTxx3iA61a78LkdpfW5NS/iDQm3qancACD1LIDCMkpZzez/ecgi9Tjz+TJSQPB
+c1MSxfXyhK6WAGTnJDh4eVSUTKCoJ/yBxb36VJNgw5gT89uPZ+IFYa1Zi7Zvnm8
fMdvs5tbn1kG3okg0Tbr77Tj4xNVcThWROUVAlF3QhA4G9FTFkzxLsf7eqoIEicT
PnnGOni36yVEGc7b0xJMjMJXQKIdqEcwgovoBEv+8HIqMJEYfihmMuWX11wnDoP7
XE6WZcKX6DaOtPASWa+GP9xVlfgpNgoo9/mcq/8roIRKUX4rK0A1m1OTzlFz2a02
ckYVi/pEZzgCo1/PPH/wrjQr9eGAic4jGwUcLc4zuoTyoLsl59WEK0eKmmheE8GJ
pw2MiZs++6B7SPcj3pf/8mIuT+P4JtLL0lpapjlv6WAQaoyioZEzdbuRG0xTuLXA
XQAIMkngK5DmJ1dodmntPq9/VXiOWWKkabclZIl+bfTTY8oDYo7cfWqT7EUKkj7p
/gd8X3f64lZ55gWz7v98AKFbSinoYHrmqZkh+2Yo+X/ILEV/eDx2bvxWs8hOEHbR
PXiO/btMgGUiT1Xg9xK3GG2NjE6UlKeUjXzuGFuN914mbXxTtagepV+D5yZg/bgv
xwTvQ/V778fgvFpeEj8PJBYRtqXaQgAvQKNBj5fKUjgcvgF/fVlx929BNqwHz14Z
BwnzJv8quwaubpS7fq8/t7SNifNniC7aB3aZNbQSdvYTnrRXLssi+7cuotIqDplD
xReHKyhBnlgSdci8tXJFzFVEfRpAq7q1NvBJ4sc24Asd8O+7X/TqLqfvykY+ymbp
R18+czuSnjJwyd6zAPMV43f4lYWtMWl3bhNsOfSCtVt+5D/ubCcT1POTMQ5F1Nm3
z/qBytQTVPw+P82w+8Sc0gbwOekhMr+vYqR2/765Cn1ChCBsnfiOvXpchv8plNsZ
3+UOQ5METypLnqEdZLDSpLmltcC3gwsi7HilnqlarTJyI58IuawdlY2lvHFMa7OJ
7T/rTVFBmefrouYmDhR5oS1mfyS9QeMXUruawiWoXo+jjOQ8XhhXR+UeRzQwvqBL
Q2JE51aKssjDC4sVaSIQ9iEucHpKGEtvt8dKN6V10SetBw8s9GwieLeIomzXWyH6
hjhJeEpZQ5tN9yMr5SP64LqgRVdjZGN9Ok7gfte9Nz9MG2LcxAIOiolvNq3d+5e3
KNYI3bc9ZUpZcGIe4QV3SUgDpoon6+p1XyClzojy/wuuEx2+geEczknAiuk04tQ8
MHXmxvjEyfGJgXY/p5xq0hSDmjImpCHrMj97kOT/xK9Xspm0x2nh2o5Q5V6sXGDb
+AZ1Fg4JdgGNkUkFWSD1gN8bmCgOtfs49UE54nk5htZrXN197IxIY/ZkhpKgVtt6
KJzqoNyZDFsosbHfTnM4LJ5kC3l7f1bB/enMXqoz0F7DLPoBjHtK20z5ERuFBcWi
g2bpgIJUTlitUFnqKN5PcZqSLcDSqrbcYF62pcwVQefpXu83MJrkN48pu+O+GKP9
Bd3xhDkOOt2N2aCd/GbBYQit8yXBE5UpHCXY/E1A/AgMOtczUhhvxATt5Ot6xk/q
zj+HMBjUT0clJnB2fUJ9O2TovdoS9pte8tN+Vd4Yx9jer8K/QIgcxDpKP0voYu38
xLtUkwxx74nXFZwABFJYfW/uqz/FNDk+Zo/teBpd0W4DOwkbKCqGGIR+3mkcJ3DD
ZmwrZMPelMFfVvnCPOMv+wjYQxq1Ic4fvjQr0ylmkcocrg2D6IjFwbeScZgPtlYT
dVMiArT4/F23vX2hXVpq57xUGU1Ylm46gZX/JXSuii0h5tGPMGGxKPBM4tgiLBG0
7Zl8rvi27JIFYSM9VXOnykgbb9f2QJWFESnMbB4WV2K/vYBLjf7uhrSIyQxARvj2
uXtD7Q8O5wFziYOMPPiutDRDUkj9sAkCI0s8rifWufeVay8VtD5pjXoyLgGPorNJ
7niPbAXgCnQtmzOgeClAXGUn1Lr9FCh4g8Zg/FvK8afyW99iUnQ1nZ5zZ62MiUnO
YgZcIP7k4JxPKkGgKOkOQfhWnCe9QcfW5ZR1Uoc8uwJpcRMllW5Fd8XoPJtsGF9f
gEQY2m6uIz54u0El6zwaNvLsdaoV0hfdCG/lFIlPMycvUAM7avKC+CsjUZudmeTe
eQyjyhOMpbCzfS+gAAD3WQxvdh5GcIiL8XWt5165JAe9IvQ5/RBwUkF9HvRqra07
TDON/4C/CuvlVLHMoLWybk2s10sEYv5zhJWH+Jscvv0mkQdciHvM8vt7mtt3+AOl
05zjgOSD0hcbFQ5vM1SzLoTnLMVuvRro6I/xTwy+ZZPMVlIlgZ8yf0gxpbWVk3pM
WbJO9zXhcoIJsIeuFSEs5hHUnJ0HPu6sw2nwC1Q01LiolDhGJKmCR+QSR1UJTduL
0KHMuytCk3V4LXNq0JLNG/hJYxcrlK505gXwzxvCsEJf+wKGriZ+VOrItMWIQqhr
6810jNPlTgtfaOxsPGvTm2nG/gkjXSW/qPwu+n2L/i4XftwiCtuEmNf3N8qEcWrh
9Lf8/b39rKgp4KtaswKtVFRG6mj9rM6rkPpCymVylZTUsWhca7TyqIefXeSr+Dca
jYL3JBXGjv+093rxkAqKxW9tX8YQ9/tU0n9j7XPkNy/a9l3OImpUaNeqOuDpmVPi
/OSvl8xPngAvYNNK0EjYjCisL81UkOl5yJ+oRUskroOBAr7QmXgYc/mJcy1bnPS9
Flv6SC0XDvJZ6XmNvztlFs9G/uw8qd2zMA6ywEL9xVu0WmwZDzdAIkr6NJ1QljKw
dEhHcjyMGv7LuKAgftO6WAE090TDQnSo6hBB1R1xK2hB8N+qwPkq55X6oKCn9XkY
Ceo2kMiUSH/OfnxgjrPS0DJ41AcODFVGAoDv149K6D5EGZ3iz7jOTqsBYAtBkN0/
C3rddeQYiHAA5xNyKT6a0OHDQvxRsmHRXUCdF/L/w7AjRLbLJk2JqyoQARYoX/pr
pBVNOR7+AGi8tCp7JwqM/TlMIyGrHxlojp5zwd2I5T6imyznc77df4F2EHc6uFkN
lTJzuEy19aNz78JxMTEJZEMkZ1JL7PRGO3aq2CduSPR7np4BAjBPMXKAX8Qqtf6n
pUL7uLyGfBvo1LiHOInt0ukQKkFZ/4l9I+KRFkKOv7nBmVtTLCqh6dCL3/u39H3G
2bFJDJUd673OwErxnJ3aLxx6Lmb627CX2TbYsh1/bVWWUD4VYTTRaY+DhDUn9slf
zZjPsITWU5P5D2AnS/6Q9iW2ZTKXV0zFvUh5JL+g/sHcllaUz5ul9Og921xR6uMi
xfHRqjzYcy1rALN0iZ/SKygpgNalR8D4MaxPxD2OxOdwUxoQ9bgUizxTH70mbavs
Yu+WCb0Tf3GoESCIK0wPtg3WLWG+fxCG4XndhjVb3FeJGdnhqlFx5nbVbstLjhq8
HJ8YvI0x1RRiOMdrwkgrbm/IXdJBlV3LtrSlBFFb3LxZoOLjgNOo3fIJ6Fs3zCIc
KR7RBnoG7sx/PYiWDKXXfPr8QN0U/luohoJY0IQvZ5kRqit9bpyaLbPP2bUkK5FT
x1ccxsT90LUVKa8OCMjdh0iK9LKVKu2+FG4i0kQeWG7FP9yHBqKqQBRdIFFkMd9U
CPDTIvkexANVfhGGjghg2aDoGiMrOJcU7ShJ81DsVScgpMybptrKrPmz3rJuKtJ2
6je6FGpPvdtDeAJFB2ZhY6YM0V72bMxuXHPWtHVBeqOvpFuW2VLU6CuMzD/A1mcE
cyjTrvr3lx8XqualwGDXA0Ldmb0NwGWTcecfG1s6TFZyEkO8g9kBmqnysteLgkTP
cCM/gvvzEOaj2e28cUx4t/qASCUhKshu7VzyMlXFQvD54CLaFpJH9FB+iJXKlz9W
WOtAHjvD5r/eCZqzLsbkZbIEmMjVXeR9RvWEVTEetlXNBSH4/955CsYBdvr//KBw
ufJfQHg3obogukQuAjJLLrQ3E5ItA0dpVfmxFVg8zmQ/jJXDkSA3tPpTAFInso9f
bLV9sm7/7F/TVMFAVzv6Nx3duGmvpc/kSxRpGy7TtetFyi6VXriLRvPSrNflQemI
bYuLRiaxj22NUR2MTujqJcNdSEZvwsha4AoD03MZpm9lqdfQzaoNCNQkacu69KEv
VXCTIBuYtjGQ6dON8tsM3NBoDCmCMuC4p4XiFwrAS54vZnI6KbMgg01RnRICe/yb
tgupSEzHUdbtPgJop/Dw2khZ/tsMSY3wbwtj6WmbRRZRJ/dHyCaE3qZdFqyLzR0n
zGUtZ+ColH9ioDtA3LwdZ6e2dECCyQMMSxPoOpXt/y506H0afpREH0Z1JP/uc1Mr
Eb+JC6fsBoya/MlsCm2Ayp86HuQ5anDaZGxPsAnZnH8xMOQ/+NLJIB9J6rXar66q
j2ZnpE/QVadduETR8kytsvzY+y8gXZgwoKp26+xE560uSAJ/weSJwR3aln6YjOc3
qkxWufijGagZ8tpLQfxYbW+/hM36TOs+0e0URW4DgUut6gAnD4vgiIpnjAj6YHKA
U8O25J+0llHoHkxhoxW/elVnD9T+gpVPoj1qcUtvbCYYQJ3Ni3T6sJp2v8HQGqBz
58I8wn6+NvV3HQ1+lhWCteRK+ocFTALHCV/bT3ZzV1O1Ed33FcwFV3Nyz6n3pE06
Duxh7U07gMWwtFBdcvGFvKBw6tCaCW9ExjGI757h5oHVnzN7OsQiYbvK4Aiz5DJO
gb5FIiRiU5lC8IUzwBsjQ19gIjGiJuNZSrFfcG/0wxRkeDxuWxYWF5LsXVXGc205
Kgp7dx9RtrtrTdGGyhxuz9au/CbGC/yQKMfJRKfOOmNtcnAx8UkOg0HfuqnpKaud
MgH3e/4c7ZSOmUr7dcah8Ny4bKDqMpH/W3PdGjpo0q/OHSQtt8gN0mVZ73IFEleU
I+LuKd8J2iksFl3Rsnq9Nh70THvwVIZxT27/lJXSBICr4eqQm33lSMDIKcQAF2r8
BnOtcp3VDNvPZZBvhKCnCMEqDTfxyNwbzuCB8DGKwSOjX5jnj7fVRbphOe+/6/Xx
BOSZ5TlxaDM1SUboTj1PrTwhtqpER8PC6F2A+hqFOI2oDPs7pTxhESoj6JfjohBn
b5oKTpUtmvcz5LLPBsiwCL5Y2EFdcXU9pdwOs9EPbpyXR/pAuRJ0RvhQ0UHq4ys1
I76OhMsDUVKIaRklgVIcF4BJcRA9/L8h0KzlZb8X2uAiS3n9WYb22z5tkwc7qckL
5XVxeJaotqWUdbMUkste9PfhntYV8M3vVL7nJytQBbstLy70DpmRpa9UKyqv+3/H
TM9eJhCC3U9l6wrupSI0WjzDXg0UN6qE9WVKNG3nHnpqwT6SBVAceafzGjl+xAhg
p/jfj/IKmPYBsmkPluiaoHtH9JQvbEiMYLPrPilIutQvFQZI77fhVZiMcVjxTn58
jEg/CHYdF5R+xoQ5wVZ3cAa3GEk53SSmWmmJNeVS5FhZa+vamI0KxW0TaodRCV7U
wTf8Zg2IgFrWddvQFHUorAanbFdzDBCZqm+m5i2uR+VC/96d2J/S9mnZUlgad4iT
DEqkETTYG6VXYwsBzWWJsZwCqRtV03mcxJu2EPw3yZzsEvGOhyVgyXr8t2T8nnz5
NQkVGLz+qLG+0s8Y9fyCDx0Cd/z6BAAkoi5kcqgA2pP1L9mMJO+x2ScN2GSuw26A
hQ/nW1jBoN+aZb8Q2VuIBcVlxAFtY7PdbQFdWDYW76UCOzrfNe+Yic4n/ycdW7rM
it4/UiFmpIZ/Cs30xMn0HLElCvFfucf+XqSOqY8oUUgoQrTEf3uf2r1fxhnvmogF
ykahTDN0C/SmAI8ZjNxE0TjuHB2tlJZYzHhc5RcasPGApinhhD3VXlQXhW9T/KiW
0Q6sz3YEvUpwyxkl3TZK5YOGIHLRjgyECaz8y152jFn4p4E2T0xmnFnNOP1NBQBz
iwtx6+rXlK4f55hcjn1lwY6Fg6/EdD/Uhq1IvSJY7HSorkEsTZgiawwekE/60s/I
3hFG0jkIyJK7UFTlOYVXvdDX/c3OlcixBryY7G83NFAK+ge4Y3zZmsAMMjwBAXNd
a63L4GqyFmPJs1FHQgaasAPbXZaJABeI8+sMZnZ0n8Y/da+kzbvngZ5Mfz/MrR/p
09m6ctWqrFexm30svwshcBTPkU8ycBE3OhqgTtg2QH7+qVjWc62bN5bG1MTT+tYl
OSIo5oJCcvjOL0Sb+kPBeU0cZzEOI/4VSnxflgb+NaiPsdZ12eF+gO93uDZsu0IS
4aP1+dNGZfm+gpyghRRhQMflL8ewINVqokIrzWqbQxbHGWUPoW535/FZicLisM4x
28HLqRTgKwBQvuGC4OvUUQEvqCs1dzNDZOuZ0kCwk0/5COaH8dPSbvbexC6cP0Lm
yhH7SJTsij4XTerVhe39jO8zlUmJ2F0y0cvZMl+fBqeYum0hc91IE2EcEjO8kk9a
6EUkHNYT1I4zzcNBNNGd6JFieDAJ/04XEbMj2Ak644iJipO0b2TmKMEm3rpE8KzC
A8fmkFDw9CCQppC1dslFA+Tp48B9CFRG///oaw5w8cYkpnaF4X7pT0T8+MrIxHaP
Ml/lm0W/ciLm1t4ApnOKnvnLQod2PLxrekvrffnw/AyOvr4vjzxlpmFH+HkI9rVO
TMYqSaDGFEb5KRr8jhPYIM0BtwuS6O/b/U2B9hn7CsHcxdl3cRk9GW8ns5+uKCTU
mPOhpdsNu8laYPX5XgE9+NF9mfaBYn0Ig3crQFQhUhcDy4B4B0DB82asfaK3xIli
WEKGETYOTj4Kq7Tt6qrsIANVNTy1BsrwxY2u6gSsWu9YFvweaVoGrwbqa1osYTuo
TOq4GlDEZ50uPPe7NoZXddZMBiblmSDPHx4snpKg8gUDs90Cln003ht/rDZXb36n
b3BILORXtkOkUU7/9sdREQ8juhoCpHgtROjzLfk4qWHW7YEcs3KLiCM0ukE9GuY7
K83yyudGCoU2VAi3aG9CrS/VPSVmT4h3K+a+O9zTIhH6nfSrwHKF/WvVQiq+AI8i
OPq7UJf2vGDw4YuOJRQWPYK+ZdE2OJDb8XzUMkVR8Ri2eC0bmdrnFk2yWS7m71e5
1U38x5E6q/5EwMqXstPAAqN2ARz1U1pB3+/4HTZ7r/z990KSQcjZPG1uNxQPgYqq
/68s64fPahHgUsQox/qEkOPHZSyjXMiu4vhKY45/O1gMAep4VyfdEPAjb3fQVAsU
4FQmVglh+Fv8Lt7OLLHXShsaXVT2ufODWuP3c6kV+UDk5ntSZDcdtXZfcj2GfZfP
/uHliqjALy+3pGDXH//Vx2w0H4FmVkwbz3/4gyHYUCN48KfZtbvV6OmqXm9x/nZu
P/CwUxKkZxEUqZEpNVFAfsa/1utoYcrJSQ8MQyirl0AHwReaa1/vVSaEkEMTRC/b
C7cIn++4g23KQzBob6tHeQg3BkXgV9E7mfG46O4egFavok9kEvYUHkzQr6vLdXIO
IMzsdbv/cFfwrbQXoeJZNkrrVTFGes49MCwQX0dk0sYMaNLibF6+353jEvAmvQtO
GjQ9PdBWaymtvzUp2MOyJJOjpg95q+Uuw7FSeOWqvN2dK6OobABDcw/b3dasNdJm
7FgfT/SLkhEfugSgA8iOhWhYTlEytZUq8tS02gpLlMcvmPOoMADLYN8Snxlo6Kgz
fvd72e9X8HA8JhimT3YiAsCMSBcHhUQdvJYYVlMmvwRNU4SED3MB9KwjWAou9e0u
vEUoI4D8bfz+nDYJTbhb9HyBUSJ3OeEFAmlejrzEIAXNJUxS5udVX4Wgj1d6qwjG
ZSUyTieyIXhGCcq4Iy9tiAswpSC/t2aW63yYkmVfMFOmllnEwq2Q76pv5C3/qCpw
UcE0+T8Ad9QPltWvmrPN4vg5m2WWiJow+BqK58o6OXiLkusL4p0GOMWNizuDtWkY
T8r0NehE3A52jt1TVNFNkKBzgepUmL8bxRj71po2at9SZ+fkHqFDmES2aNGBvbNt
so0gzDu8YnZezHKzfN0Xlmq5fjtsUeppK/1FwZArwinlx+ManyiFUvfNZD3Zpd1M
Lz9kSNs1gIaF+XDD8RiBTpcSI6wxN9X2ON2Os00Wev/oSFkDZYqkPqX8GQNtxslH
e+w0tVeILEBYFqPEgCuRWOIuNp8Dt+3YXfRZHuqWi6kjh9sq4eadOoUAnC/nVUPd
AudCY39BvOrDqkMqhLDo668z9ntJ5/EoGhTNdbwFXoonsSkXyfhxUG7nhdzsQpvT
1fv0qVZlKg+Iwl6WOQSj8W0PeSYqaM/dB3/vrPF2TgsdMCQlGgy53h0JD9eyFDu/
SfH4VNfrhiY2bJqgAfw5ejdMhveCm2fWSBasHZevzSPA4gm/c9yhxgQvWwQ5ltYD
O3es1kYLhlbkosrggWQgXuMs/4NHe3H4RU70qE7n/VOotq3NsUmB301VYLe47AZ+
Ldw9+9bbCLKfHFHCmeigtapPN5puVLLmfgnMIKAV1V/twmwJ5DAqfLq3y8a+NVUz
HRrp8PqHjgbCa1nePq6V6dBnV48W3u8MYK1xHLq/qhwtsa3087K/iXxLkGpFl0lK
JF4JOoJKTLsWiHeBuocfABQPzciZPqVG7sXkVTNJealoDuw9Chwew12jJhFRsc29
wcxpyxzXAHXued7goZ05F8gVkVXATPLxFfx+WUJY2y26xGyFlKQCYyP4dm3G2uuD
FcS47XByl7OsyafR46ayfm0o1auV92AD9nTgKIShVmqzkqs/l2oPmARHnV5n/5Sh
98ADnwaz2zkvxnJas0stqweaycXfEUdGReaQZecderq7gKTBEgfcB+LdnbAsZMue
N6RiImTCEi5wy6IM8XffT1tCiSacyy9Rsx13K0vnofuEK9EkpO6QZCRNqSxO25lm
hEIvsINNolQXO52IilZFSxdahXaGSz4xNdZIZJpc0dsKdNyYJnDG8bLl4Oi8MxEs
IIZIcsIF5B8x3baIDAqScwMA9U8ySa6CekCo7qs/q6NkJ3lwvHrRufmpq63/CE5U
eIEjOko4pLDf4AE8NTlTUcH0daYGpWzZRWusa4/oesCYlqKVN2PoMUiIl/8xaPDp
Lvcw0tDF59tWl3qgOQSyVSp80NEPjPXaifNNfWNzlNNNsAJyn0pp4lFq4MgnDjiW
two2cYfDTg1pkosj6+me3CdksHKfwQ9m/w3NRvIM+CIvsdrC7VMyPua9GgeMQqnt
8TXxpnR4qIzYx8PWrdDcpuYK2twyioiJKEMLHftsLHvDDk4YKZX1o4VmIiIgRTDO
qDvoT9KnVtKTpoUP+oIiM+WqCyLJxWA+JmBmG1vtsIS5PXPBl945gGCTG96iCFD5
xdgCnOulEhKPU3ZPj9doGKbm/XXzOHLME33oz2kWNCNAAolOLlDi7tZDZYpTcPIn
/yIaLdyQRdv58LuYlc36PHEG1uSY4zNYwboh7FdA7FnaCBAOLzMAmfgA9DQDtEDh
Gee96OLNJZxCUNPyQKVJPcKMpPVvik/KqpprHUmBRPDmoQ/8iS26iNdAXF0L/yMt
L9zONGbkFcFmOEtCjMXYTtxkOsRizAyd2A73v5ig306BH9xzyeJ/fl4jeuSiUN3w
sPb8M/W7KhP58jrrsnuOdPvN32vvR60kbyZMUl5FmkyevlChu88p+NfVIopQhBdJ
CLd0zpK6AGcJXlij5CsooEz5LQ3GTzNZbF3R1ugwcZ3wzyFu/YIm1Wpf8gEhV+LJ
AF8gVBlX24vB9FYzRMEcCxYvkYhT+aDzEmPDvV0s2QRV5wj7U9F0FylbvAzdA+vw
fs9lWepWteP0wLpDU7f+9Cubj+FTaYQTTP8k8CTEYF8L0z1bTTnvlA4NM/MnvUI9
DduLwJ16gYo44b7KvRUyVajolZ5loVv9fNyyz8SYwLp4qyOjI+ChekKSqfKpMdcw
lNKGhpFZ9Z1QGq7Vq4+D4r2KMmL1ln1SSW7NnfTeIny3nzwCKn8lxXEGsFM+ZpcD
nxaJhoOaR1UyKk3SzoKqtuw93RbsIWlWywMOFrnzF1riFIj50TZTSviaUxu4e17m
DkST2NHYFk6wyXBwAhDssgqYCfgbpL87vmd+q4AF2HsTTWjuNyuRUr8WfiJlqsuG
OqItmmxP6FI3rFu2oMonZW3Lae9l5Pmzs5AOBzC2j0vSodQa5v5FcpE0GnjflPxe
PPSBxwpYT2U80YWx0VutaoET4viSiyH8E/vL9cVD1JDd689235Nz4HCPQEqHidgI
MTNe3GmWhsVYZHaIj0T4SOQTJsHR5Veuy0B/2oGkuFrWPHqREqj1hXpduZbpwqOU
gSow1xhkKXbfWShuzaek9DXRPTAftwT+ZLYjYmaHwWk/tgAl6y3CfSod609E55Q1
J+uTiDQ5JwQs92nOr2+azdnbCx6KY5TXGg5HltY07s3QsFyZYT71C/+NwdG5+K+p
Sg9D+qZa1GQeHrLnKY7G0MMEd+qUJMboHoJNQaTwohOxXRnoST87ppORSgUTQlW7
3KmUCt77Ad7T48Syds5y499exp1C36dhGlHFmp9wR2786CkcjqH2izRt8TyFmpMt
jFR2DUqpSu19PvRIxppf32+4SqH7nPYxHuUfiRL0ubrbvYhJCKJxUjnQISf3a5qz
5X34rBK9Tmjv+pP+Q5xSIW77dZHxv9EhbAbxCAmU5hme6R0himsf6OF0Whk5flus
M3j8QDcWYDPfQ0GQq6M240FkPQenS52ymxKJjs0j7lsO8Zdpb4tbTEy+/qIOLbT6
IXYik1iwpz/aT5PspUOVYvE0ICtFAkyZiPe2H7t5XBcpWfEkTte3bca4trEOj+KX
npiQqa0Rra/ZFa0s/jk71w0xVHrDWVyw6sADWUQi6i7+35HcK7jrcriaA0B5W56w
BS9hnsnaNz6S5Ckb/svA8+Cya8jGcDIL7ST8Jg3SOgxcTDY8OCJ05ugxIew49q5v
gsDsbmkoTacGuXAHLgiKy3+evmHWPS9aDU9bic9Fg4VezfH8CwgI420NJH9esqhd
J3lDXiZdiefOiaAsYb19df9TdwJ89O3o8UPrHJQJYREyseC2ZqykEAh0gP7fzVEf
JmVAXVwXQkZv0zO5lc4FSPOKzxDX6+dYZlkKeTedo2iIG9W66Y4ZvnKpG+ErMKvp
UIyvjiFmdWur8jPlKXVNz03r81leRte7ZJZekKRiMC29g9IYwZwrsYAzcx9km55k
M8vUjvPk0zhnkBDyl9mxf/lcSHlULxN+aJoVIClGcnj4AnLbvQjz5FTwQapJ63S4
sQsDXsJFAgS1vC3uWwjYO7GDnMtnrRGTUzbeP8grK02dNDBb3JBHcpK4oYn7PE37
M6I2DFyOqsSEnJmRvp/EGHKzY4ua9sr9hi7sDzCtWtW1KvJ6cx34qn60dvCnmT9K
0O2HqU6nzuSrEJ3mSGVzGBzww7AuRdS3k3DkAPRlBqdwy5xn3uE52m4OMzq5safl
/QoZ4dDzQ5RQKpxKP33CxnE3AEr/m15dUGFHKeGBWpc+wUYMQCN5TwyljP5G3ymp
CogExQZDRVkFLcwBsAkUbwXHh1I1cARXtKhAcOFjzAyF5l73JpMa5baZpQcV+IGE
qIfAmTYO/puagggwo76jp+3t1IFfzZDHDOWQ+88DbTixnIfIsv/0itLO+mBasuZh
nmAixJr4YWCphFTDvRgFR22Zw8RFd995J7QR4LkHXKHQRfSA1E+WN7tRbIW650mN
5jgHuYU9FM9/K/wf8fv+i+hbgixtzpSkE5byijjt/ncn24+GPvrwbpEn4DnNS9VR
hOK+GZR2nuoZtlXPIzs5AeUzAQJV6sp42OsR4DLqC5yehwwhLYD6FVGIl7El4aAi
8RRfJyXF2vVMoV0kpHafH/0nj8w9St+29bE2yJL8eCyAEcOBYI57zDSfJ7bF0Yy2
bEOzbWVC/wXV0VrdxTnYgyrxgsRvRWEt6ZdB5B5rddWtzlGL4XX9e44JGVQ0qGtt
UCoyDkgjjg/69IcxK6/XkqVYo8jr9OkxYcf8kgK2v/nm6HvCVUUFrrqGm+7LERT0
ey3xjXByywVvs1RSoh2iK/5TWM+cOxa5+fJFWZFEfqNvzf//oeOHylV0dpqYIAoT
g9SoOAJBEgdwNuyOAtf2Z87qE8yVOvH0kLKqkajYkmH8t8KeMRudEPWdjjlc/F2b
pKiFaMM8ZJTG6Vw1Dws9HXzIYgOg8Mj4FilXbH2NpXxQSc/G/j+r1Af9wFle7GY3
6p9GGFCjHz8nTGjNvpzVTnnZy04svmMAW7m3TDGVoLLaUiwmb/pC/SxmTnRGtWdx
bzAoF+/yjCfqylyM+rqr1s2oSJKsGbF5IjjE2xvr3Tn0dcOPHw4dTuHqnIUkb7hF
cjaoyCa5XK01fsfcSkFiAhFhpNYpkAEbP2wrDxiCLg90qBrmteKPh+FtWY1D+D3y
LfGMa8vHva+8Ay94kVSMgMAKB4hH/LO6ZKMmASrnoFcQnudTN+gTLkFkFnbCdlvo
3krB+7/E9ieBFiSOb7NV1B1p/jnN8Mi6SndcNQt0QrQxXzDExrvAGvVWhvUrKhV6
Q57mm+UKpfiqDtAb+Ks9+RWt5yUeRHYWj3SaImxwXlppiBjjLT4CBsjVMCQxRvXH
ebxD5g/3VmVr/rNSI5SXavjR/Js+3kd4hq4S6oT34Z9IHLCIRsEAJFhMl/K4YcYY
IuMC5R8JSJHIPEOaksqPxDE6mPWLZxfXkT3/bXECioHE5hNPg8H9CcQ6aFUonRR4
Lh7QVHAI0l5vE1ueg8FJNSnidyCHqTLRJitvMCL+yEspCV/12NcM2RGs42tpPJ+w
vmygxMEDsKjwMIE7ILtEbG6huwSbTY2F4cckzA0ArA2ddKwGJCN6jUqk4U7W6N57
CuUPPOerss8N0KLRjycrcw30AJkwdqI8yrn8Y4H0Sk8oT/iuDxeHBsZyiMwyM773
7nK5yJD1W6FPx/i9lelEcQKnceaX9xLlnqLCe92LoWObdaXhsNLj3o7YkTeMiY2l
HXdolHgWN5tFKLUkSMHGnK84uYdojElDWCSL6u6nZJoP/WCXB+0OxI+Msrp1hBhO
J3/mmIOXFX+xk9i9o2sdqfMNneSBZ2PB9sYyJ3aSVsf3YXN6c1HPgL5jo1yxcjdZ
B7mtEyHZN9EtXgfsRwkb3Xxv/anjmqvlaZgFHi74BvjkQXFFZwVtLYoxqhcD/zfu
17SaWc7fEelBLEHrY98VEcOAGJTyDj1U4HHldPwt1SidMDqdbSmJ7Fny1Pcwk/od
KyazdCuG3BbsVplyMvR907bO1RbpgC0HXZjgZ+pFMBiogrngozKrprGmya86jLU+
bp/EwrcvmFnJ2g7LhVVu2/U5tSiOkcMTM4kSAu0wzRXXI5nx31ca37+LcmQyHZgS
Ytl+cY14mx2dSJNunkZSfgaOnqUtos6dgvw4HRczxz9zQW40ZXikhpZmTaM1/Pxn
K/eAjc8SuRLet0C2O4O9eWvNHjf4HpsoWMWEAuuGnBONUTeg+ffksKkq5z9/jkTc
vuF8Aq1jq4GsOpU+/hJ5/osSD1PXT664h+1N0Wu0HgoaOeV/ADDQ7kmoutBIElyq
P13ysCdYMk5zMtKC7cjqzrNhhn9/XcZG4lTtw5WNwYz05bzRrvUKC0RwAPEBcRGi
YwV8gG+djVMbKQF7UwTPU+KHj3+abSryRnTvbuOAGZQ4ah88JteS3yWKwJ8sdsLo
Av9ul0QCpVQQBfl4Cbuk+aPkb6H7Uy2EZlOUiHMRUon7QQSZIRm8d2nUu4/w1DS9
RfZJcb3pT56mOPhiMchOzC8fBn5hYk562vPi11v9Wo7ecPBvNN+YCscx2IrSFmBr
ualmQEjf7WvOUhoasLy+fQ4k2B/9YIgnJJGg+Nk5XknDh5ClVsmXiDUwkUgLwS0H
x8B8CWrxkS+DSYYRlekTIySjP0OH5dLYpJIRm0vOR0CPlF8quZnlXlEXlv2127jM
JBb/63lL49nnCSCBsCX8OymGRdA933pamgxHY3k+n8g8zmb8JE3ZhZxirH6SNn5V
finJEVw8KwcEw2bQAErP/812XBKxTS/i5C7vMoO0/loYu+C0ZJxETvqtmNHZaJMQ
bMeZRYX0tYzTQ6x3wL5FrFN9thKTjdARfcs8HHiUzehi4mcrmOjIa+tHRNyDXUQZ
A/psmBL6oewmukaoFMASO842E11XRc/WOmrJAp601v9t58JJZ+opXt/kvVljo/I/
/uVtRcZJHQoGz2U9yhjm/1r/ngo7nc4pKeRhcMr8ct0bz+1yiOJVWToJxMGKZXkK
hgE9XnWIIV2wcMagH9u7XFzbz4X9EBxCajMoLsGI/ZK8ZihU6IX2qX2tO1kPqvC3
KdzvsmNJqCGgQfPKoZJTWb8+JUII9SIQCoqPEIss+Wx9oYxY04e6WW6wIlIYoS3t
+7E9K6fDBFIQ7XALe0FJxjzNuLJ2tq12Wi+eQbDMzOChBDWZe/P/Dr03XU4uUtvf
EiKuYWXqVIkQLbzhiNkZ7gCVJXqnBw4TLbwUz1MIV95a5cYD4YGc6WAjrK9lJ036
HI0R/y83L0x3wsT3ht2Diz77ezotNNBvdbx8GvcLbSmwMaBoBPyr1Omzmrrt+qKE
1n223wItzwvKNkKAeyBqU5jylhKEUO5xQ4hyvUaoG18oDIpQMRv9U44VXUabAOnC
HxqXE9X/DD197V5OThMcjlONHLaK1QtJQg6ld7OEZ38Ss3QgsYLoB5ebzsnB+p7x
rBYyBYH7df5RvfueykApFK+DTJyaeOKxqIFStSQpWYKjEeZsD4gNuvQ30YFYR3x6
33SQgMSJ/JcLKdcEB3CW1T0F8GM9mikn4jiyHJFbHnjazDxVFmVdhqSzZ0AhS04S
yortXk+oJ17slxO4uEdLGeggb2W+M5BOroDm2FkLIHVo8E6gryn2UGMW9AEHEaF8
CKJSOJ2oilvruebviP8Tjsl1UOThWw+xrnwKede8BVtSnajFvOlh+s4qf9kbqcsj
2wDhBPfj7dtrPYbIvbkFxpW6VbFK1+qogLWfFl9T7ETbhKvUsOxVbc+RtltDiTzf
bB/+y0GGPzlRVJ1QuFtB6ADIFyqr2j6F9e/U7kjuYwGaAESsAjHCotJluWwAAk1M
xnVxGjphwYNqAn0mrwG0QWnIbQQRilNBOQIugNcx2GRZMk1kFtvO3RY2DKPbVJT6
wgIuVzx+jYzubGYERlyj+CK/mGpjQvyrWh4w/ITHmCEimwXmo5mchoA06CqyqowN
qD3wolb7/06iO2sSEEbg/Z2BRgan3cYlC6B4lIxXXhHqpf3oYfOCragzPPwpUBmH
6YuXC/M5I1BRXuaT0YnBglqbU5NUrUqpOjv0ywi0Gz60J4J8uMhkhzQKYW1ouGZh
Xz2Geq2tG3PSKk2p0P/qQ1tWr6lFKDOoqkle7pTHCacdOVmhNhLbE1il8si8ryNJ
G8X6T5Wg38AjhC0WdqggPo/Df+jua+GbbJtqOovEZHIm/UycPQkzPunBNbzSQgpe
tlwIjBpsH9k+0l3YtCwaZlFdfFe91Tfw/sx7xFBF07sXTQxy6kIQFuES2AUUMqQ+
N+R3i4tli4xr5RQ8GvMoTB5Yhlusd5fv4RfSTtONZpkIHkcNJ+D6CdmRLLMk4zKO
OhsSMXd964VPZffyaCLlQI09pW/ZsG4E3EJaw6SCq0dl+ck1RhLq/rJC5mK6f5c3
sHYrxtMfU78x85VltBNzsiHUY8dBSpyWPFEBYOcHNNst/9W5/VNSxSs66L5Cn4K7
b/yos0fPld3DepWw96ax73e1PXYIuQkemNEgGrSeeaDl0teovQRjZz+uX1dsUAYn
CmVL939kwmC4hhv7S0cSzWaDkN7JLAwhzYnKoCLirNubwOD955kv0vSuHmAsgq3v
X3wukWUG1ZHNWal4gfrnoUL9HxLDpraW0ID5CmyXUWSDJK96oPBKXolDQzg0f5aC
S/XJCSFH4jbELETDfozDJCH6Uj0M1oCfEK6czW0kaitbEBjWXspexQilr0qdrbkF
vqu0f8GxvwTP8bf875p6Gj5aqg3xx3Hl1lIS1hpMgy91ywi0HxJvYEfwlIU/85SD
SPnNKjSrnffFBWZAsuThAUfyn7oH1B7a7gQQKnXKiMXFVrNFLIWutLvAqDAQcC5Z
6OPddN1p2BIA9nsdByTgm8YrjsV+9pdq/2jr/rwCntv8R3T2YphICSZUoZSFdxUY
QlvXMbRSRClLVrBXop72uTb01kZbqvqcsRmoj2z2f8cPIknqGTiAyZ+MXuXUaKMT
iY7HEySm7ilIpmJZdw5lG3ikinbwlBe3yqtw7SVYZnhRUQZphdh+F7STVqSTEtlD
9O4NBcUHmzq7P5AXrA0uADioQz8ShB8QNKU3iK9X/opqw18bH7dNVUhJ0PjJR1xV
YQtk8Zoo8wlncDVmuD/Be5+3S9wNoeOkzqHcWt0TPO3mOcQVjiCI1rlNvoYEzUaS
LNUPSQT2VMgO5M/QLI5mm1OUY0FduzD6tzKC8ImUpmPWno0jcUuSrl0DVvI7SqG+
G7O3HiNbvH8qk2cg3/0oEngXb1oHVnnWETTbFKH0o2665+Ldkx99AMzs4OncKgEV
xtflmd9mpeEKNgDPx9Ccqtw/2qHpsna1L66esO5sZ0tHJUIQxh0kNDCe24ca68As
OTtr+yMkwpSDct9OavKwwmW7mlRQOHOL250KuGpxp/xiT5/JybhlYh9nORpRTirX
bolfzGdDqBy3RVVkxCJjTymRevzXSlYo5JDlsy2kbMLSqdww/JCZ8SL0ko4ImjEr
e9NM/Iix/b1m4kocc3XRU5EKKAcWJYdKPKqeHIjOdz4ET64Hkn3mREkQWTcXL0tl
dbWUO0V1muqLAew7C2vA5dWf6dWhgvoqXLZjF5vHhGAi5+F1rzPTSPBpxvoFZOM0
fiMsXP0S8vxf4+fFYeywCsHhqVRaEPtO/TO+u/qrPxx6lmHxC/ePJS9b3YXOkK0E
ZCAW9tW3GjXtjwoZPdPvNhx9zyRkNYp5Vmbed9RO5H7MuQuBI59epydjDyce7XE7
wcFx4GfKI7nzK29VOcX7B43GsBN/bWqUdBrSqC2Gzs4RgiNHTkv6xzUp8UHWNXrQ
QEXF+2vdQOi+VDzPdfbwmLjm0Psg9gEHmMsHfGoN+lwLX+QpZPLfHPfgWnRRJdAV
QutQolWDnHCAPgY/Xo9fK9Z410dO0xUNEij3foUA2dgWDj9TGRseRQrEQ1LmBOvI
PabWYrBk6lmXijWSbiT3qOlIu/lyTz5jRuX9MHDYms+jRhiw1ttsdiC2bJE15dc1
vCQyEYvi22LY1aFaY67RReliVE7SJgGxnzla90Y+o/Ki7dHdjKnnwc/KcVw1XSAN
nWif2d+fBhqRSJDODNXZRB6HxXxFFaKb6k69I/xOE3HxaE7TOhEj2gFccihYhRpg
sV1kaB0ZedGEtB9w63qPRZVhVA0szEIHTsjN2MtWJsIPBiqFCs/llqgs8mxpkYyd
q3j5czRFYeJME4VSNC7tH3gST8X/QTte3X5pMmVpWNsEeUNEjivC3BF36EitA2+l
EV1I1LFV/c+ABuuPYUyfxes8mByd6QoPXCzX74d76Qy/sicehsa/OJJk7Y6qKUM1
TwrF5pE2S8OY8tbSdcJynS52LWlqqVP5rfvlT4CGl0VWzcO4n1VcfDK74VUcuP7l
9C6R8dIKEEBgRoQqt92D2zDpxYhnuDF8fQq59+qjS9JN4YJdu5JC1wKSaQxKupYA
wplHt5e4ua9pda2XbAoRFc6pa6y4TjugIRhazo2sT+ljQvg32vMF+fs99ZBlcJWT
TidbNRaA0ewRQDDIsUraIARqWIhTiDu15ZXz+WoY7C8+I59XDCSEEOJJV2TX83L3
QnVMV7DLHnmPjO05O3mXqJAzT+tsLaEb/i78rhuaLCmpg8mSPSUN26i1WK5ydzw5
qxG3ivnZjlxikCLVYxyTsrBITn5SgCFwNRlRtIKl4bNbVmHxDLcjFnOW7LYHu3e0
aIxh1A14AwZZbjSFMPfIxc/Js7DMthktZb36ZryLksgP7YmzglvyD4pg5AtBQt7s
KQP7ujbNL7Qf8LMI0AlOHq+KmxYG82xwFhc9nuVxidhIKYT1Q78WZ+01JEgCSvUC
IUvnToOEQL8Fs0i7t/UE6bQnjRtCltdq9BTQwZ0Gc3tMakP6MC0rZm9ptzMBslQI
AflAExODEeOFlPLp04OAuy37oJ7KEJwJ97LZSYwj7lu0tC+8WN5k0iwVEtTMdxIo
C29K6ay4Vn5rXnwh3+EpJ+FOQzE2UnKPzabkE9Liz60FrDUwge9xVRyyIkQu9tGw
xgusLepF5DhazNtu9kJjq9sR4yhfZE+UYRDNfS2mp9Fdaf62koUh4Pdd/owhi27Y
KR5FDMgWrKyZfIVhd1ooK/Y2lnc3flp0W9ynWu9EQt4EFtmewftOeVAoaRg9tCXr
ERePt5iRhko2+aSYcMgBKP0osE9PA1yz4dzrE/ZDqqplFqkZITcnUR58aS9thNAM
hOIgT3+Rf6E495C+1AvwLo3kJTuwq6TgUejh4j5kHxACySr2VujUR5YPE6bt3UjE
7B+aOrfIXe2qwOfCoavehNNtLCMPJY62ow1V48lvVY2gx9OHuWjA+naiRDU3HqZI
WjBYEpYbnuNtp8wev+t0dvM0aB2yHC8YbyLsvpcqRarSxtAOlxIt6wO/P1xOfCU4
5DWdvxoefZBVrgywnhMJrCcIN4+3ADXsxX2rLog3PbODcmUqriLq+KHErZ9EIi/l
RkGe+HqTkkACHDIUiwlPv1Kv3FDMJXUWbbvLorDem0l3QAqtWyhX3XFZNVJvPYqI
/wAZN+mx5mGLYgWdNMv/eLO/ZuxCw0by0JYen1M7c8Px1JTxLCvpIK5SXd06B0Rx
HcJHMadr73siwkfQh2G9KXlHYIB49xUVqkwBxu68w7Fp8UBAAZu87FYiUHIBLpqk
goB7nJySPv8T/Ym+kwj0jqyG5VklGdjl8j1hP0XpeA/shG2N6krFjEAne6gLmjk+
0YOViOyRLp6Wn/81H8+ag4G1WJKJJ3s3H7zdp7n3jURDKx84c8s5JFkTlbpcAttv
NSkTfESrhqyXqgoBVw4KnJPLCCuXzq2vHR65LSXAPDn8OxLxzB3j6AFlzfVvU5rf
IfWrgfmrpZ0PK2o1Xue2xs6wYRyZgBwDJlDz+r1QOol6zSiF0LFRldT/6IhcJl/s
60SL8CJurY+RJ0Puv6yzUgtMunS2eV8sbrS8UN307OB+G6CgpkCUnQrDFjQlR+GH
auxvmsLDaoQm9gCkpmaPZ4bNrgveSwzMbQekDH4CKYm8XMEiyOcNVzOskgVifo8F
L7zSTk62Lsq7wTS7plYWhHs3TkckBUIsGFH6/KgVuzxUObdLsiClrtelDnnper+J
kzIlvcCyqYA9jBoaQesOx1TRJCtcgUzzKEmZADAWVaxA+SB4zd4NRsWb3I3YLxpF
wZo4klbsLyenwakqKvrAB4Z0i5h0yZ5Iql+FmSWtKsBWD6YzbH52FpcBgxbNFzOV
6cmMm4mAE4qS4eZ10PiU21Kjqu4t/fjvv464hGZWSS4ZQOVaM8iRjC885+Xd4GMu
yNQurEw1b2Y+wmGk3LdRa2BTyXmwHjVfGELNR7kvFgCFBLAZOVeQpi71uuojBJyv
6HmReXUlhxwA0BX9W+i9gwFDDNGr/yNRiz+6cKTPzb5X+X4ym4+z+RN1lPCuc81V
oPj724JRnLQVraFINS3IZaGIQmqdN04aMslKma0SoP/Uc+QFPxhNIfGJpshkV7Vw
D+A2huw75EkAbl6VfvGG8JPuHFgf/nsRQMuAzgq5u1Ex5apkL/5HF7EWNJLYk0JD
MEqbJa7mQZHkKvm0X8Egi3VbdlamHyO7qapDBMCLlq1F4tX6GynnGzJ6XFir65ca
BebVtOtM+HAMQo8AEeOPklWpcfS6+qZjorDEgxHL7MJ4pu47RmHvCK+tIqWamo1V
lq4gILGgojTzlmPUK8OlY2LaWqc1rrgWtaHaNkdxWsl5YrpAEFKwE6r1rtSBb0Xh
FjQQkQtrCl+HiCdy1PiVSIC3l9uge/x2C+eakDgVzJOVzwerqaAJQfwkQuWVrxQH
lEbp33YTVZRLtkWU+SwFwzApNnklofO3Z7cuuVNQlTCLFjqBbdV9ft1KxD8HmLs/
FIMI8/KvN80gV/aWOahUeHXN/DkhDEiSUmX5j0jCJ2Ga5EE4NFrCKhsGFxZR4m5H
+c+ZmiclQOHC+cYFPzZuYgJyR/dGz71tZfhKNbbi2Exw6FHRaFTCgs4mn8g6ZmqC
XNy3fZtOELf2xZKA9zzlGgQXIzvJSs7gjrSm6kWXRtxQ6joLXXgzSREkn04RTKBT
t8yP3hUOn+H68S+MDWkxjv3p5j7gwx9HCw/5OEHxSec9NweuC/sbvSs68kRohVFX
/tdrGXpqhD3pzUf7QyAuF96fgZhD6jGvxvYTdzqstugvmNJTbIGi1N4IqvaU4dak
5GbXq/VSk+rJmqi+d/c0LSnrkFHcWQf8D+VHC50/Zts4Y30YZMcBe+eFKCRtVbwG
qoUhOLica7RJ1Is2lk9t4WRCnKsr55Ix9mzAjd9+QiVIyiu41KrXOePg62uugD8e
zWYILroOmXbZ1SevXVIoQ6uuZj7I7dShOBmCRxch5WXfxvMDlqEzO5ipD+y3s5d1
Xz44wWUvtiuFP/BmB/pqU9Mli+T0g0bhkUpj8dFeuiGiecmfRSe70e9wPIb9KV+i
r6Q1Uj/+18VlpcWGJgGaiHSYz3f4cMt33oAvsOAftkL4n4nfu8p51DDU6X/2q9ME
t8UtOJMR5NK1xKedwoudJ4jXv2wpZWXYd99a9C0Qjl0FhZ+vBJvo2mxuCMk3Y/wC
VFrD4mqC4hEaHTXnpUno15unG1nO5I8bHjAkeHZVihcpzzxHNxONT+UbZ+MG85gw
zQ49CFW7gags2n5xfpW+mcwgOHT9GqNdP2u8eGjSHmro2Av2L1WTO6aRNqBQqFSg
ea7bn+ZbimqtUwUDt64IEyTt2ty4BgL3XUQw9r2O+4Kvwg1ZDN98hHz/twFUsCQ/
oIeggBmZKmb08I3ysLBSOh9HKETF9lVsKh4tkmpxChjYRmGZ1okcpOdxtdtLryfI
Lb6xVnNK+Hs2r0PIkTR/4uyfEcy0iI+bHWIjxd2ohjhNAKQZS/aq50mghuKObQYz
qnZqScS28Yy7c8bcIVatzG3ZmutQgBJ46Jx0ertNZTFOjpHOqwOSNWimK8EoEPb5
76hOU1P0frAvZmjA482Q12lMflvERaanG+yzgBXphjLvDU0MG/uL7kEWNf1bfIYt
Z5IFOcQV8HFEVzRk6Pkwgf18MiB2NblCMf87D5CU4ccjVPbC5QsBwdF8G9d+fLSE
kmn9E36RD76EyEReTHQeuhNHOfMc60QBgT5vUZDF1wF7yfJYVBjtg00MAUG/nN64
3lzqcPAOuB5XlRCZxqLaXYM51wdQWSfsOwmAWRjCKs63gQeAec8kXXU1GI/hLhrB
QZXaowWKX9WK5NfTXd3aP2+1cX2K+suEkHE00s3BRSRgayOsNSELV14FvLk6SiJG
U7ewHBiTC3J12ib0eHIlUFBp0iB11oc8wHSA7GU/pI5p3MMR0qdJGLxjdmC8qPF3
Zy59Jn19UOewPyblvY+QpmuT+S26TJBd3F/cgikhsTFMrW+xXr2V6cXRg9DUZ3Z5
55JZ8JqrLWngnLQuKn/kAyjwj9l4lWY6a3HuooPpb4fVNQbNwChEwiuAX6nhkoiO
EJN7K95DQeIrHdcL3YFnrK5FhHUdis1FeAlbNW/XpEdw+730xwv/XbauSvPKryAm
NaaS1EAMKlWvOaELUJV40M6KndH75d6iNmWwmdLJEVd1Y6551vK+uQIL6gSo6ja8
I17iGSbCeWULKUIWinsciUJOJTc/9WZiTuZs7ia9W5Q2W/lNtT9cPkdQmXdsf2Rf
PC1Z9YuYWotewiBgHpx9EAmXJj4h/Lfctq2evphMDMc1acNZOhONNCDb8RsUGsZY
HoMavJkyPOe/5r0DVrPjOu8rpuHUvCW1BenHBWl2jSYVxN4j54B2RqPCJgQAEwED
CGmNnacpG/ZPdYEdYYzWDhPCQiEB5KJL9ExH+eXBGnCiTGTWwmAfG+6hC7pol7+n
609rkCHNGGSj3tXfaD45EWYSwpGxQwYLhx+mcBvRxx+QwTmj9iHaC/78MlQheig1
G4Eft/9rXZveijwi8nmnFFeHnobZTIDZk2YTcYohzj12wqHCcihGSet4+YV4u5d9
WyUsA9erAvf3Q8mQSsJjP2/pa1xokH53LWnMDiVCt8t5COYPsHEtOruU1S4sfyP0
ZKr8uD4HKmsrGOczyjyNhRDX53ybnhtA5kPCvyRRBM+HOfjwc+KZWiDYbQsYyrUZ
vQKhj7P4WGrtLXcRW9JueBRt3C8D4Eap+B5ZfHkNTwgNlHpZJXCFYLdzEr9VARnM
RKpAjZ7MFZ1RqeNnih89kvm0MsAHpZC96lKSMFcczY0dP9Af2AuQ665z2b2jDZWP
1hKPX3vmfHICkiX3EhpKXywxi4kWoS1fl/eaxe+/uMhY7oEt0VLTdQw8NTVdolLn
bGlC6f+qae66gzVmdP1hP3o9yzdFBNKOXpIQvuEH6RyPZkFoTuqTLXSSWRtF/yYD
/PaQAhz8GhiokjYr6cI7hGTr4XTryRNOiJArpHj+OKjGa9qTmCssx6q+8roFJBtC
72F4oyiXtXI54VYnlVT0LfCrGOo7sMokAE6o+1XFyAbaDZabuWqh/3UT/DdR9SOq
uiXR8Cw/b8jgOHwTMrCkrgPWHWhWefmegGdhsEZ2fv5hgah2JPSGglud+tF7ZsNV
b6nDG6mKO1QmV5JsWDr1qLUUUKIp3CWXf7+G1GABQLynse8fnkFnu8124B1aLPWy
i4biTAAyZ5bcbRLumsV4J+JFBecpOCn1Z2AQ7YoJqcry6I/LIuaEls4xGrG83Dn+
/MJMAbGAnjrq+wgEAMhE9s+/RWm4fdoL8Ba4LDzKK1bfBrUNYntcmCrc9d5FEyoz
Tt/gQQIZGZ5HK/WNT3/WRapN8UVaQoEx4wjUYUyiKCCpPioaf5dJDTDKliL4Ed4p
oElM7DDf5PHkhByUPS+JDfAuEFBDBc/Xv6DEYLikFMPag+FKLh0FYxGG4rp9xELe
OcQJ5rWZN0FVfAXVsDbzF0A5sHtlo9heMRifnv9NBhUcKxt3ybEbD7VB2aCqb25p
EGu1NExpobdHBLgi+ymaQzIMUNBDvkkABvP1/4jUwG8dfKalo/J5/uLs0QoHgsc/
/MeVCsWy1oTKVBZG8izvzxM4vPKvEDBQEYSnTWYXK2moTOfzU8V9c3Z+YC3bGVL6
1TT95iXxA3LkH0RJuTzEspL0rcBHl9/NXza7rrLmZ5E2D3+mwsPYeq5dMwsoYqUe
YHJevvysQ5LouCPzq8ZuT42qq2RbGJNOuun7AHyFpqwDfvi+3mo9O8yOabRK9FUT
1SyRBY5LJGi/+Fnrou0sB0JOLpKBbhJRleXTnotBU6UDfe6KGrjoLeNtp82xTcZP
226lDJaNqCtRT0ZBRa9QYY9s9Cj2I4QGQpCaQX1PoeBZ2ovfVcPvyOf9RllME/71
L9hJVEK03biT3E/m0JHAShG7t09ht0/NDo/CUkVg56DtMxkcQ/HbYyq0rmuBrG7h
esa6Bsdj8+VfZjOzvKAhOhD4Pc6Qfd1CBRGw/XY4vIpfasYYdlkVzPCwCW1Plv3t
tQn1j4wm1xa9rNtg4/qew+FK3STkYHHaGhLeDZR9Y53A8MHbwub2kRqEf0T95Z8E
82KncHh9CKO7RFImTtew3Fe+InzoBqhUWL6IZEC17vwoBvehm6OGnpij2u+mzXVv
ISywvWMJ4lmx47QqhYrlaJmIfrCD3eKrXivAGrD2WYyMCkwhGVZzsj4Y36o5umq6
OsvBqbeT79AjDqMmCFCOXwuLEZQSTKi2nqFZLXObajLOoZJYBQK86M25a0K11Dfv
Bi/NBpju8L9fTZU37vvFj3FeE3TXI9ayWHlOb8r4uTpZGNc6afECOY9fk2cU4Ln+
iWtRtbwbqLaE3CKuwJSVNQ7n72Jz4dKuGxvDP2h9bPQ4ax8b929Ti3KQFhJGxtLn
vjP1YP/wARwxT2bWTTaH8LbJ80OV0+7ZJAa8JdghDBqXp439IR4zbTEbCsa+1OJl
TMH/vJuHMwjCwLDH1MxLENp1JP711rLFt+VB3h2SXwaeQ8fAGG/YdXyJ5X5yQruS
/errGogyQKXBc3QLxEN6y/c0wXaoZN126n8AxPGfzfiKvlT0Q9t7bYH/XGGTXJRR
CEb2ZmOCXMr+Pj0v5cAKkKs3FXx1UypPNOywOR9zM20JcjpwLAKKE3B3d2H6yyRm
dvpK6fkTdwMuFdPTG85PPLB1UngZK6ixaRCPf5UcH0y4hDiLICsyPL2eTFGuMCOr
rXGuZpFPBdeK04XxyE26N/+hNpRL26cJ+a1RXEfBe9VCxfnzBz7lo2udx+8K5262
y9MPF5RCQQD7i1GIu7E/OKyIzOnt4DOOD08Ct4KdPKFu/vrmODQ2VbBk/tmpPFwQ
r9emnNZxQgxtQxKPMM+WX+D1Ykph+wspNnplnez7EtRebvsI3HcEdmSotOxgOjpP
5DhVPvIrwrTa10Jf8BsKsd62GVzmXrOCqaTfVIw47MFnEpS8rhp2Fqm8CjiEfFwe
bL4R3r34GQJZhGJOsgpnMWP30yhxapsOYZ3FD3/OeVXxIea4Y6fcB7xD+DR5XP50
8gjXAujp3Kqp81Y37MPN8oIkGUyyXcNKsFsxizWXfx+EAfAvv3oIfunsp9LC5OwZ
M6nxedvif2eF2HG6sBmeFi/dse/iJM4yWxHgwca3Ub2eNw27JiKp491VgveI/TSe
joRgvCU/CWCsDHGwe1BhQn0fQohX9GNmbQ3f8QpYEhLAaPgiD+6CPKwBnv59FCYW
xYV7qq1pvTTKGzst5xLjOEA4Hv41G+IgigRGDVMqk2s/ZYMbtRy+/UqcK5zIrbOA
nbx/asQ8M30h/l88RvoY6uzQm5BnAI3jUOboczTaWj7WIbIxuuhj5Siu+d9bsJFz
B1pgbFML5Ducyk3y24adAmzWRpHUmLu6xGY+OQ/+wua5c/eSG1tXgxaE0qJ6FFqE
dMOV8pBaHwbLDoqYazU4avaDE4bWlq9wu/BPnHpxwvP/w/rQqdDCcuREPOwDjISS
+8Q1MuH0xixiV3iEcOZoCHmy8OQLLue5K3gOnNLQGIdsC96gTyYDMS33vj+bVFwR
tqeQ+WEmxIEchFCPTxju5GE1LDAhT/zdNMhjglJGtQpTrtwcI6ESCGJlxW/LeAPL
1+eYuc+Hsng5iIQPmVvrLqjwBijCeD+R2TkruWKV0vG9tao95dQsCm+NSuW4C/la
7dNWnk6sIigBCCQ+uHC6DJtFPyn8lq2kYe9scKKzb9E8NZQnViXci03HBXJywyOf
Lebuky8WntFZE/2HWVW26pTJoz33myGYWiOWKOaZIMMUL3jGOU5i4C2xfZPLSOTM
6n8oFZWL+sgSf52rzLAcGLBS9L2jtWeKfKX9PPirk+aSh9nZ8lgdtfwu3XfvS2Bu
osfEf3rWUI2v2iW4Oid7pxNICbI6hzoKr5KTnb8O79+2FdnYKSQBZGm/pVmh0HVq
Yxyf7KYvfG9XHdiGQmIp2Rdw/o9t9tm/mG0BqMN1Src0TqE6WfO7jZ4e1btaLije
J1HAqxfLZyPDX1hj7T9PB+XUzYeBwlNpZGYAZ9cC2TcoE6Lh9n5gqbBv6XE/S1vG
8O3cWfIza/Ub0hh90pOYewpVh6tt4k3pljj1JyxfAIcwyQzxg7Ka+DV77oALW1PP
popB0YoiTciSwFQ6dLDazjKPvMcXZgq5+IxvvXX/xEYVXefZCbIOoeGiOLNTr6ul
j9pCuiQq/kE1ALVBobgkCLyn+dOMsHqeMp+knPuGuIVSJI0oZb/HTlp8123bEF/O
QV6+C3Imnkp0DM9d4TxZOPjVHqIt6idd+gkYMf4xUhR/G1o9zqTjDOWtp60Rpvsd
ySxQmqgbLE/bYPsqa95L3OANKRWBHKX8ML+V4TohXYTVwHcFbcdLmX6JOIgMTMiK
go1V2pTrpe02YqlaCcfWwnVpUCge//hl49Hq0teVp+3SnUnKBw01Gcec5hjsUj+J
o41qW+qcElhSLMFbN7Dc8pmmPWpGc2niyBoaBM3zZ6RS6RK0zU0pazKeaRSKH7lD
uohbqd/QXUtsAWaXgpfrCON2Uuuido+iitW8fNUx8IljD6aF56lNqqBQmg5+W/54
Ubip3qiPTzXbaYuAUmAc0Bd2OLo7RhQtg3Wjwku/0D5zq+0WsZSJINrsrpxXIoQS
Yo55Qx8fGBgIV7v53gvqYK2DtkUMil4qs7jsaHgx8/RbA4CdGI43CIjrCvvW9YxD
eHrxYnOXO28qPAFQYEqKKhpBDd8OtcmpKpvQGX1IN7tRUxYmICOu3FBNSc5GuXY9
PEl4gB0fNeRKzBsX1Ix9DUAVTfhn0XLMpcY3s2TY+AMF8/MJA/4ECsPmIdFuI2yu
/jcLLxej+noAThfADJlOpe9gfdyEX852KXsgVRPtK07Wry2Epvef5bscy5LTw+y3
GtDMF64k/vkzITUVh8sd1IyysuIg73vJJrktHPbBR0zGdeahd2s2sY1OfpFJ11iT
aCdW9S02scwia2N7Homga6khtpIEtylhHfKt9NBGJAE799nwiS5MUg7azdZ6gfCP
Uwjq7lL5cNCXvDofTOjG19ULrBCI2BlepGrGlCOPaIpbROzZz+QhfGtYDnxmS25f
H40sAbHvQfRAcmIiNYiVfkASQ5Owkj2j04lvfJUki3uzkgMmfA7Qmi/RB4R9HSs/
bRFDzjWdFhnVdx9mJ4jDhwhHdm77pShRMDTlSiBPOZG/L+LUaC3Zz1whCVPId+Bi
j5AlHng11UNEbQGEuV0iDri6C/27UuC+RL9klytzHj4wO0G5J1VqdfW0Sr007tlZ
huczyzLBssG49aAxnJA38PkKL40Nrd2NoESIFoXsBDvT98/TgwG3pPi3Eej/GJPc
xkh8QwtJx26F2GtsqwDCb6nREMCQsRA6hrZ3hC+OO0tfwWQuPs6OddysK0t9m/7G
JF1siDEVznyZLvHwlyc9QQ7GU4LqEV1YoxyimXhXpbef8Ee60l4OUfa7YYqY99Bi
6Ky2cujMOAvS2CKx416iGGZsQWZGj9X0wa2dEQ/Or0PqUHTl3VajIm1jr39x3/86
PWXAvIW3K2WlNwLJrx4DkyL+cx5UNksjQInoPUo9Z/HSftngFf2/IbIul2ZvCvcV
LMgrCQxrEsPYPPPz/xx+a4/hRhOUPs7Jd6CBQxyy9qpslBbCycYMzr9425WCEkB/
BkbxJdA30emX5Zi4yd8sKCJjQ5IkC+cM0iED50CfeGu5C3Js4oPJjFkgg/1DGyxA
ctvD2g+DnWUjpqiV4JacJlI1v51Z+MS0f56QbybtGihdL+bws3jsE17fCkmpFXDr
59AsPZp+lvFle5ducgMtuDyJ7IaOQ3MbwLYjuka3VOUPx+VsVz+GsBJHXd/MI/EB
BdlWJrW/qP5L4+wGqEogJ0hptOb3ka2r4yikhZBOILGID4EB7x9P7cXmu8FAc2d9
McHnoHTMvagN5TwitdEG/8Q8YRSqg0SUdP5Yhx4hJ4LZ6KNFu25DyAhGhJPolvxH
vuxOs+JF3b3FlEtp/ZFMDglDcRFBQBALUqAycJ0oHWf6IjfnkgpsaDCxDTTF4Nmh
+WCcT6xkooyC3XKj8bBBGKvOygHm/4L/ZzWS++WdCPf/9TnviOjLjy0TSOu+/nO+
5pXkGW7q3la+CVaE14hWF7KD+t5Slu8G5xkWsu7rLPnQYSnWu5Z0lyDMKz8wN7Pz
5MlzH8JR+W/E0KPd22AyGr/kIXMha/72XtDdjiDHFbMB1AZ05YmNTCw1OZw+kv+a
GctELZxcLcbUKBgWf3qf5iCXIAy/dT7a/U1rEBE5lpLI0wJJMq8bn9hTGCNkXXjo
wNXBRGcVeeoGEIqEiv2GNaZ5Mecz6po5Nbx3qMssWz3oy3Tg8+lUwHE+nnNfHoRT
6TTtaXrrAtW6S3rK905CZhsbPzQGElmNtebxAi6y0ENxM97h6KxcXbJebFazPZaf
IezpZ4zQK2+AWa5ujM12xW6IIZQzcXsyb8F5NrqtINmhqccGu7DHiipmn5pjoSI/
Gt4vho+O00TLB6bOE5uziDsCfq6gRc9p9uNAa7kri97MZ273QJKbhvTYr6xhiU/P
Qoa8tSKrC4pxFPWcdJuAzaL92W/EtUsFyt/jyu1j9EYIQ3FpGElYmu63AiFhTfj2
ppHPNYwanVdU7B+Ea5fIjBIOkE5wKyryrb+e/HoSy98rR64ox80QKLgpd9qSY6EV
BJi+g9XBrEBk6HVeEXktHOFqXPIAvpAsOuX+7/HcmEmMdnpcp7TadM6ZV8KLn7Q+
tt/xR6EG7UQzpS77hIennz9A5zhRpvSlEY74XuPvBbWO6cOgnhiDU2aEoZGiuY7g
R0qOTx26cwF+sVoiAPfJH9JxsG0OQ2gxTvNi5wOWPttCaFB1zrHcfSd7HbCU9XIE
XoUWrdfqLfnO90eB3R3s35eHH9mwbPfN+pDx49tW1BMKcbUTNsNzRdhR2CXUSmRX
UjA4YOix6zrUuEO5IX7rbEYsjnOa/hrqASdBsg4JqXvB+ELyKiayB9n2UXuF3emL
TeddvdSBh3+48St9VHonZag4iThNPzTX4QnktO/BnVo13jrb0NG8HM5xLrgILfEP
Jkt0hE7ycrardZV4FTIEQjZXk1P9vmOhl+qLF75iQh106j6ty1RkN6fWqLfghG2s
YmXYTnoIHcUH1SMuP8hmGQMBgZ+AtVMfgLsm+uSCEzEl2ysZ7MotfoUdBfOU5PPd
likCAsjvhnPfWM5PQIpdcQqjR3kKEfT6wXTldHbtf87Nw8X67iWdAV5kU45EkRne
+MwwWVSUITfgAteNUKSiUVsYsIvarLU4lXiaG1DYgZq7k2/fYkC5mr9C/Bwe/k+/
ihhi3oT7upEykhJp1WZEGR8UmE9LbUycevXLOjYg1UvWn8pCtSoIgYfPHATkWEZn
pTfq43dWPdaXoxErp94Oc4IOPRYnCVsCBKK8kCAEwfwmU9rB8CWnJZbtN0vgUTK4
jOpuN0uzvdEiKlo5JGJ/M9wlShWCZ2q3BQKd0cVW6D9FZguRnvwAOzTPeeHwEens
uGLOi4nzcH4v+TVccB8DU9bwuDIim58WSnaZ/ClhAwMU+D5oNNRwSjZDO9sY9NZd
z1kaMqdVmCFOlawp1ajy00xR8dt0jNzeOQH9u4SP/ATXRNfW0E9dKL194aFOWti+
T23oHyZL4ooQn4v1A6crBNzGZVnfztug6HAxM7EEu0yuiE8tA6h3FpP1/pdq7Xj/
oOG8J60/anSClZ/VTrkSpME/cJS+25QXkmiGCnFu7P2z2QIl0EGlf4mpP3gRDQSz
r/Fo1IOezA4iDIv95voH/9OLTmec3RJGeJwoi3xt4iYwoI51UciAgsXWByK7rJRz
BRpahIZX4oDP6AspSmiHeG3yayNSuhsWtxLiJw6UCi5z0MRQXD+ngCv05vXYnbKN
iA/qOZIK+LBmohR/7tbvWB2p0Ycf9HpPqXaIpJBp8vXIqZ1zpVtFEES40uBvN3Vk
tGaBgnRf+/e5vrI1d6LAnBivODDTOBCL07iMh/Eqr5fvxs9i10w0j+IBztl6xyr+
86ClQ+H9UABwW/hiozNNBwXwyesj5D+S5IQtLh5eStOX7bAuFptXMyliZ77aWSZ8
euTdVI8CoBzBOlrtOtQWiKfvCsma3UKedg6jK85PEtlc7y1d2QvKKMx92zpeFs5j
NhE0tHjwKBfmG2oROesbRkAbvBmXgwZ0scQ2rqSYw2DZGauWVwm0SoTIhBJP2Re7
qeHK7QTDihs3yR66mCD6wvAvgZI7sQplt8LEGfKv7yDo4hN3Xg9Lmcnn9fdoBqxB
XkVgH9qiCRZ9kjteoQ2IlJIOMKQgnYFPQ7tK03yAPW7510OZz11zYxqnpEUwaCt0
5R3gqsQ5RWl6jSQiwS1xQ977EFIrd4oCMvC1B3Sd8HMi5xd7wmpAwrXQkAy3KPCX
pe1luU3y1VhCsIRs85H7tRNQ0QOCpWzUL+K9JZVH1KJLvBOy27tGaO8c9OpC4ShG
89nGjKos/R+EPvOeoFj2Y26fHjKRTLxFdTpGyvlOJHWrBWqoAPesWge1TBxAhFKg
l3XZ2SyttewLSJJQEcCpNrCcWjKQFlJ3neV4kicxiDNEFSXWrZIntHQWFtUg18ih
BCF0E+h89pcdxfUentPWV/wznXYgHz3OyDRoRtx8HJwLOw+1E6IJMw2iXkz6Uf49
/vRUaY9FFSzcG0Ve2wk+U8FP7gdkw8TqnCaHbhUg3kq68PWl4T92VWnSQkXU6cGu
AcnKz0026aAgrHSNM3PLvQOBdR6NU4l3HheHhHf1xBh3lXONmtDMOXn6osAPaVzK
5YE5GPOOfoBzEiVf7DgTJBNPH/7Xf98MoncdzNwLkOxEmQtHUZPcXfiKdHC1f77g
RxgB6w86y+gBvl5wBJuVNHHaDn6bZBWcwFg8bqfmaadrT31K6fKvhYAWWSyNPbZa
hM9+sjc4ca+aLl97QSJwtmqfgv7f8sevdRz2b0WosukoOCSqdQxlRN1CqVFRF9uK
/KGm9k76KC+DPBCKcPUgTzP9d5wVib3bwPPZsuduLqb+sEnqx+UtNCg9068/e+oz
QwIVsib8g2A1txnd8Q7BL71HvmQKz+QWC0NlFE5IGo8A2n8kjJWTzvppLV7C+WjZ
uP+/Lai2NdXAHhL2mV9mh9IVkW0K5W/ULRwJxGYOtz/R5xd99DgEwPBu52i8Koz6
VG08njJs3pV5NvDQVAljVny6DjjanbP7szSmtd4WunYq2i0tMv5hXEcgyo7z5aXf
0IkAfkBSENQ2gpGbo5CaG2Gh9/NSqBv4ZPzkqXPwxONTDh4FLG2NapwS6r1TqR70
ziNlQqbyiIkJRs4z7LSlNEmanFQvSCiBvq5HuC8gV4fumx6tf8IMkZdXpDRqwNFU
utPlrmjMjYxysImEudqOft7vGfibH1Adj/sZeoBD9pOxGZ0ijeSnyFBhHGTXhNia
h/IjsWowPNhoWxdnUVeAUo4ehku+wQyJp0UmdwOyMFKhYSZRGgI4Ml8C25mNXpno
GtPVnI1WAe4a0TPGp6fYObY7pLEoxO0fy6/ZbT+IXmyK9U9h1TaXMTkamoGSKqel
vDZxcjTv2DJuDqKsrZLy0540/P/qELUAuL1x6jF++Md1HuATr6pFL/1F2C6rhHEW
BCNsO8UGj9l32Wzq5T30DcPoc01fa7bbOQ2uO+88AwS4R5KyCimvDi9avRLF/jI3
3PxWqVl+/SRlUIlSya1e/K7eVKrUQRd1jS8haA5uTr6cP0djZ7ux4g4vuIOJNgTm
UgcUilI7S8oCDYQLTkTjSdZXFC12e2jJkwAHrroGfeDaa0a/Z35SJAYopzepTbG0
JWn5Tu2AyJdVnywcJ7vCILXeFdsupjPh8INXMtPRzDystG7WQccWuD1ClcHQHWT6
bU8mFxKGRv8CKnYjguwY9V1WDPJUpSCO7BlXA589di1KJGVDcc+OtnW+DPetcoMo
xTzhxLwkwwo6FEZ/C776zOsp8ZualJ9rSj2Digs1HgOkcagcjvPXck+gFzn5E2sv
U63Cj/PXK/nti16wjaMV01qpoNhwiOqBvY5o/a2b45jXDBZxeWtAbBLSaoW+DZKq
QQpGlsXH1kQmy1f5bmY/Qw0/hQFcFKzEQwTRK0y0mfLS8TR00T5dFWzNhfcFIdMh
j/21irqeyJdtIG03iezLJp65sv9KVISU1y7w/Ph0Fl7R1aSkqFvPBbUHVaj7Jfca
i6ag3QUFieD4QFk1a3cVbuuW8uGdMbTcOQzEXAe3pmOIbnUJ43gs9innXF1RDcue
Qh0TkKKjIHBuIwbOvTIqDZFLdnhrGdPsCkkOYBX2Deh5CEOiJyVCl8xBRJApZ1A1
ZmrefJXyQ33aEAReqohX0/iQRCc6FJeoRkcdqRNM13hLtIRO7a4O4NFmQv65097y
IGkmH6uFuGAufgz14CdpDU2pJsiMywA0HHE5O0gpjVB5+ycDps2LfgvtEbTL4nXX
0ahG93NoLiYWQ3UCnwN5YOJ5LRS2wpgzeV7FEy5rWt9Jkc26VKXFg17TEUf0zPUg
PiWgT5U10sGsRFeSto9H+XNCcnGQJ2Or9xxPttW0YgmSwx0tn9MoysdOdqA6asyW
d3TtRWQWuh2cM4u1k10A+1CRpO1HCnbXYxtaoG6Gg4a6TC5kWR9Iaq0oWJq0sMVV
t77Phlu3EWzH02qQX3tl9jHZJJSfP8zW1j3O0L+SPwf8RgryTJp4MVhVAHKkT3Nm
Zx7ysQs66tYisjrLCxzuJH8x86RHgMpim9AbKYscsUM31bJTfKT+qJojzMFpbgAC
yQe7xHI9dwY1VZXN0ANhwy59X4Sia7iMCtz1fhNw1q8ETAXlPj+Lvr6jYzAtFA70
xoAMzm0DvMI4SJcpcioEORZ5YhJbK2g3bk91FeJKdHHJJeHz/HeBd2+nILe5UhbC
qdBHxXguAv3brF310oe1mTjrTwBcQZit/+yBMqe4vLOMWJagWx2AUY9iBWTfJQKh
4wHwxXqSpNYbhat8xufFvR91m17tqIzx3yfcGHpxaYORx7Gbf+dIdp5v32U7O2Vb
/yshPyEAR4vZTlKdgcd+sBlBLaQj5s6HJq82r1nhGROA+82Ax69ugv4ENkQnTuEN
z3fgWOUOtytFrFIh4vOTPpNS7xOCW+KQgMR9s9bgcn626tN2yAIG7tJv4q7tY3vt
CL26f3AokRiorW9dCfgdcVJK8wmKb+vUzdSucetHU/lBovkyXMqm1YfqMtiCqFec
yeJnWFNBtmwYWp3Ws+O7zr9doExo1yojw22n38fhc3NNw+BkI0AEh4a6pOdUO+dW
edJ/UutM76axq8di2u+x5wPcwfT0Wt9prVM66HNc+eRkr/mLkeklRtLXpg26t1++
pFnzib3d+KbUU5kpkLvdgs+cOJswPudGa0J7N7qr5l7CfH2sYNjSvYK3eLKHs3/t
3XhmKxp0zcB6GunwvEA+GyhSflojITPiezyZSsDrAMAvxL0i0WcgIGOLnI7tOdgc
MbAKQ9e+vfbBCp2PDq/7BLaUxJv+Tm45HDSR6nILjldlkR6gFvaLkMmiVQG9LBKu
NQYCcIlFfw/w5pOLROHCTXrQvNE/paDBEUh/rqCULp0/PTQAxEak5G97qPnbCVk6
HQ3AW+Z/jeCjlrKOhIagukwQFwPN9GTjYDJ8/3NpAWSCIHb54SMuddTkuXdOD/sZ
DJfSaTjdpyObI1XeMjuUDs/CWTixAZLQHTk9ok25NLwPny2st0WyzwMs1t1v6yHc
73ifq9eJqwmS+wMjkkfNKjHwMyI+Qc6EdeEtqUwvRE0kiRYQDHQV0iblCnb5Txmi
8p8F6XQYYUAaYL8lOnV1BebweVkeURkC5VshG2r9gJ2CTZW1vjpenzQ3EYTL2O7T
hExyhQiP6s/KcH7fWkSVH5AEZTgrQT2pKZB71LyRHnDHvQJGmNiBKMXw/etULBlE
qo5qQpQeX65KvwnAV2KDom9nEMUq7qs4G7az/CUpexZI5g/Vt99h4YEpuPW1mYju
5qcb6/LWLglI1AbwCdwTjApCEHWlcM+3Z0M/cCVIUFcV/giJhzl3P1Ui93RSxk80
4urR0gzD7U+CyT6TfpvtzXwP6QpvN4sGhULYOprx2j6qdX2BG0j4T4xHvxkHcXNR
+q8+iam5Da2FKhfFmOcSgKhp0mQLAknj6bcqNaO9SXW9EJnpnaNC8hCE+0c2QmBi
2197OrLO6NdnWsNvfhUOP9iFOIErzHeVND1soeyjrgdrbkzR4N9vcsxB8YEjVXOj
+6Y44hB2PeaiTJPMGi4+4hso6nFmXYpJA9jG4jNc4ebdDasOKKV/uypez8Vo90Gw
PBuVTCoFOLA6Q9fDyXIMw7aDGZRfJ+gXtSfaYl82efTuxzne/ycFkFOgGWy8tzaD
+qd192BkFhYnsGvRFYvefw42J4C76VhY632t78lmUpHvkuv70APyOiS8tzFswm3d
v0S7MQnUYNMTbnHKbXRKXUNHdOD3eWV2wagnnbGXsbzdMoBwJEdk0dr7hjN3uoPN
Ce8O1ZT8b1qltT2fzhSaljOBaFRBIqRwgJFh96VcHHT7qgzgeMVTE2WeVgCT/0AC
IGy8Rw3FDmgtakbw3cFRvR3750mdfA9vZxyMyYx2JvVOrCVpG8BcoKGuid9UpjOx
69wg829otS3t2g39T79qBWCDgfhi8dgdeOUOFm0E2ZppyuYAIqBIcLKJ9KD+p5Yz
h7Qlp/RpvfH9hDB4HD0ERFs8ci8oKaJ9EFAb5yBbvVHy0EC4uGpeYUBvnkNYzqof
z7Vear90VzfBA9tOx5LUJV3grMcmunVH8fyslSYLKAVSM1HKnS0pTi7dTZOXSwqg
lL/TCPCv+tC76XSKve2nSvV6XjSn2z3aS8I2nQ+XQSunQo+5vbG68T3+tr8b8Rva
qAzCO6nQ0432zwILvnJfeEsfWNyLDMb+HarGB86ZzjjOM2zX7s1vbE2LrcfUqfot
Saf1YmIF0UayyMp2K2BKEC3BXMXNJ0mMYXqPwk6XxZn0uif3Wh6YDpEizeGW0cvg
aP8yGpTxJPBy4Id4cFrfiIcmhXgkaFr8EoJHU2utZb/8QtCIxANDXjF4pGasg0pZ
IWFXTjU15/OKXhDGRgVelQGdPqVaWQWJ3bRVQlUvKVAh8E3f6cUbMbzYfLdzHzNZ
hpdZuat7M5CANZ1k2byMCDElftVIYaGRhy0MsahDrRmHhUABNHycFixPSsP9Y900
Lf+b5HLERndgb814nzTfNw1GY/6kSinRAKRskC6G0EDFLrHf8jsFp5X/lApTbWA5
YO9hhgvf7V1VmwASKVcqyW2LS3qV5IelkdKBaVst54jcM4ACg5DYzNc4871MCpPT
mKSY+0RB+Hky3V1x33BpjxINFfj2jW1YPM2fIo+uE3r1o8m2LtyQSbvmLUGUWc7W
+md6mmag8JKYsk8S640P5wWrEep3MrEPqa9Sbm4tK+EHVh/7Y3Lh6vmqPZ1Y8ObQ
PbtiYHztLGURYMOljEz6DnQjyZ70Gf1MafhGRJhnuercqWw4JwDApQl9skl0d2VN
APLZnSkyxH2hHNx7KIRge+3RamvdLdSKNMqulUTL7DCdK1dlZ24MEYQ+hhyrKeE+
4p6fkMaNwdABmYWcGz4gTBWDhj9nP7vjy2TLZu9sumDN1/IygsWBbkjCAVcY/U9z
rPyHgeKsy/4OZlvSI5H/VCxc3pZvAOK1F8cWzv/zMw8HWyQpvnTYUdrz4NjUREyw
zwsfxhSCywYmH7U5E/0HyZ69xT9tMkpoJLc7HC7ngt57ZTPhHFkFJebk1QZPhLWQ
a92k6LQEWB4oFP/0Yp1sGr3hXLSADp0rtkoLLUUXmP5n3pa1Td9dV5czxzVLcpDt
3lLDzZ/jyqOZpqyW4gmvMTyNcqOTXcGfdn+2xn38+jwm0wLO5Ox0wTQShdFHNfhJ
PiHHko5A1t9uLzCufmoRaLg1PHLTow7nlRg7dWjbVZ4skLKqH4jeoJbLvmCQASOh
ZsKf9Jwd5UAvGDRjxeemVsh3byQTtQ8Gh1poI8hq99aNzvkTcAvVOxYq/BzcxAjs
jMUBDjKv+BFVNoIHxr1qiYDTMN8wE5k2On5ej+1yHHFlZXNTYx3CZnt6ZYtjUjqn
xurL1C7euzbRb21q2p1JRdz/wx0deR69byhhGqnFQr5NtgFWAOH/0QzZmSYPqxSI
yqtXfiBY+2EIuTr7/iGgbJ37z3hpRo+9LxObreoC8R13y0qmG7nLsHuRO7xLAoFU
IKa0SQ1uRrt+O5Pg4pXH4WDBoDFUQB3s/mPAtR07iVuUXmJyx65u72eV3ZvOENdW
3kQQtUBlZO0z8XurPXd24alBzrOPT6YEhgn3BvlpnoZqh1S9zq0GFglgMTBEP5xG
kJ13ws5NqdO6Nv+uyq5D0Cj3qmiiKt45ezNUvIDhFensHZ8XWgGG0xXQlEawk25z
T74qgP6l58ahsczUM6q0Lo6WgxVeRyUx1yxCQfjYig38pFjbNM/41fn5rn0uHgWN
o6QW2/VZTdx1xSYPGT7eWZ96Ol7Jj5QJLK9hldIIRkWpyUOpEF7n964hxdP0zrgi
pw7VYN9QJ6IWv0DNaiUJm5gG0ozzZlbycAOsRVb7hXxmXsbpPDs+4QjlIrsMVHIc
xc6gOoOUdL01Uzmsbqt24W5c7CgMIEr77Lwx0b52PAqNo70uP7ZKrvvIX89xZMqe
xMr0BoUPdT0T9pjO7BiZxGM3P4C/GyCk7+M1aT8LdXKJjFiHlxodGN5siRdm4kZB
E4NQRfujSdPnXExzoSzYsvznZZO7Nms2MXk+0GxvtKgnZ2hSI5LxyIcKhKcF66Mj
ak8K2/sWcUA0v1JahDYhPrbxsE0X0Y+o3bIkWkzzel83oZPMuJ1mDLUQnuqjtqMn
xv+4B/uwVk0Ihpn0aD4RAAqwxElj25/OqW78ISnxrd5Kyg1H8awJOzD29CUrHR8M
7dPbkVzXnBKs0NFG1MxSRdCLPQ7LGc0B18FsbK7b++ecqxDlnj+MAtVWsCNgXJMG
2XkWooofDGQ81UA6/tQbdUc6+G2aM2q+6pejPgKn0IaYYiBUxaFqRl6fnvE+RauE
JtfQO1wGC0yzqwqrIpTTcVWSL6GUXUsFZlpLxp0Kfbb2YrIv04VanqVBCYDhvgjD
8Ve4bYpQMgVqq1NK/zem2KqISCgqtkNEIenIL3P2LPRmuETPdLwBx6SKsWF3bXFc
lZnUIKtdDRqQRnShL0rUAIt8Co3IvW8C8owVUSy6kczVakozpMtCGsMJTxHvN4Nc
o1Xc2PISVpFYWqwtjdTeW4C2IJIRMKyR3C8NpNlicw4JGHdXsA2AOPufEHTWn48g
GTBjwy9yBzt+KILltb67veFoqJKw8o6U73bD0xNpZJASUJKo/mAnzZ0nXXxU5qpt
HT4Zb89XRGr/emjMm9D2vt0MYZywcaajtAdKI3KpFLxoaJ0339flOZeeZZVAjw6D
VZ49+0rGe5LRMEyIc+aZQ1waaemk/YMSlZv4zbAL+ddLjV2f8H8gMBzaghLxegzo
zQBOnOlFnkFpL6iOE3tZppJby2+6hnoqyVgoOAHZ3iS5LcxaHnDJ8SOi9zuOPPU9
cYMY7ZqvcGwxCTr4N1Kwu+InYF1ugHLEsPC2wvVy9/BuxTs72WWFb/478CZpr/y6
gu3iVf7chkWMyBJtiNeBHIQ/DfCJwgE8un8irVjM81RqYxPevTGc9Oe5DhTQRiiL
XinQhwk9kcz2VVvBbd9DB1IrqvUnP9m+M4R9VPAulLesVy+RNqXsi6dEMKeHIrWW
B6Y0Xw8vUBBPngpv77FQRbVNUm0GX2AhxIuUKvQnqZxxDQ3pHmhcDYF46trGR5vr
xsZXY8F7hwF7WLJSVCiNQ1Pdmk2XNmzqFNkDZO4OrwCXaQN5Ha1p+4qkZc6Y/aDJ
65cOe0grJUNdnASLB1LyZzAt7njkV/rzAo+tKEyEkmNjiywih7/yCODdJOkaABBQ
nEc3zcClMmHfoTVSd7jA+7exlLPhahS1GECDpt+viGuk9dD0NiYFIdwDKBp1+LlN
eTbgLeiGUuCMsIRo65mx0nxddGQ3ltyd08PVBXKdKJSCY3YtcCRQK9yXYeRXvBTK
XB4kzfPW7AhNbr39w914LuND1xiRz5n7Z1oE5zF0MkdZl93a7Pk33GF9sqFO8Y57
5Ud6GTLiMM8iCC+U97gdN5x1sgIbwp1Hy8g6dy1ayij0AlqtsQQTFX6SfHoORwzF
klH97E/MryUzD6K1ZkXR7rFh1Jfz/VtwoaknoY7WdtM4f61xHTJXS6WdQSqsIy5H
Cg9m3SUAmX/pP8v77rIdX61odHQrjU9m9S9N+cWwa3/f5SnieqgSon1aQukXEKF8
AR00VzG+W8jqyWImJGnbbThUS9ZwnmyF6EaiXcuQjqdjgIIw5Or4AGFVuQtgUIrw
GGAcqh+p5K/KTEfAI92VZpvj8korEUruaI+GyJfqSdgcfeCNhaeo/rYrH+ri46Jl
0iEW/ZXVuTeFd+1BwMOI5c4MDRk2Pcgcc8jh2nZmExN2HH0fSNJZ/6JBwOWToTRu
gVW37/hd5qDCaovMff+V6n88+3CchEqFsSJyIXiv8I+ekfM4BzivUjkpfMsN/7pp
491+ytfjGr6EvO+JNz1eskL/qrVzrmdbeWlO8NVI5f0DK3cepIphuPx/kJ6ky+3+
nj38LsaGW4YrGHsxffmZmCGaTDG7pc1N6d1V8vivEpQrsCF0H3gDCKowgHTaSpWy
TDtPQXXwdqu1oeZSg9klrdKUnnxMPnQYR/+H3NB2BP2GkuieITorM/KWC8jizTHP
LEpSg3s2y7gRkAPao8r3+1FV7ILm74l0k75pVOEda3SH/6toqgIPLqd8bDTgObwO
n71KJWpHukLj3v483CvQo0oCIU7+zXfMuTZ79PyjChK3khmhZOe7cQo/GBS2dn2c
7ezvOHuRJhRLgkqPGBL0enQcoOLm+41nGloLuZmrOLhxqYMF/nizDDOOT4P6Y6mc
4hKhZXgCE/Lx9bnKsAhRB99yBbUfNxdqC9kWkHDMJtjP7g2MBnuuGv2hWBQ58Q4N
/MXjXUw1GfZWWa6NTFRecwkIEQG4ilmt2nF/5gypIeUW2za+RnMh8SAzMcmSEPfl
7vzmLX6EmrUUxyNjcGUCzw5gsF6jFSI2Pc9tN/ExvVMYCfS3ck/tocdJzlwgCxcJ
G+qdZF4rtgUlNXpGnCUbUUSghOYSGWj4vdBU0qD4RpgVAJlUNjsmO28ODlydCPe5
3HfZjx/7BRaikQCPvanNu4Zv4+dOZRw/MGfX1yVnGRkXAuDmu4gMndFCqmuYHce5
3PMo6sF5jLLtLp6tNVU3+nTzHMzUt6T5WTqCuaxUJREKV6Gvu0RswlDqqtU1Jt2U
kP48y3SUm4q9qUeNayZw8xF9Bi2c+kZgpiBuY/1H651XVwdsFbFArB/Dmyi6UOLC
zfCDKPFqCe9WQm35ONKClAiWdWbXbwlcBnCN4E5cAwmEbE7SqDH2WN9cn4uz8bsn
KIwShcYAfJDcMnUBMVlUjkPq+XsYRwgxYQm0p0Txxoplo2jhb/M/cI2Mpih3HF0Z
Nr9H2EV2Wss9lPN4bzMEiQqSEWWwVRrJhu1NE80+KzOiAg21hxagbiwd28Y5d5Fq
pGu3wuU136cLwT1x1Ugq4LCNjft4rJiKREmjjDZmpWtqH9nq2qOmwqtD1Mzo6YU1
rJ4OdSq1Pdw9EOUTDUP5ij3w4vU2tuCzuNokvxSJYk8/5RFowyENX99QKMA9fD5W
lORK2rtyqmL7JEb/THezKkX9wfn33IEfbPBPDLjJnJDE064WvKf7YQi198MRejRg
+51Y7AYGdVtPoNZx+tNDujd7ExOjVaFQS8ZG/FDXewVf7qxsoHRGsR2k7XsPulY2
AWH7+qqfSkhoLUkwiqQl34geTS7R+/Nppfmtb2uiGdo7u6dcjTtwWoTN4FlfNRyM
Xuur4Msj/DloQEhiBJ77jRma6f6nK5WuFJjWr8oFIBJocnG+hcSMrl0trK7OiPvu
FClEN0dpJn0COUedfhL8EzLQQHPxaIArBWgDveOmeXC5af4//t1MgJF/tljIjHRw
IrF3nXb+AVHFBs8hqgX7wwv7l0n8kHv11LPJZVxngM3TrFvwgi4COwZGHPhkj6VC
I8je+3NTSS+DEPkrZSCfds8ZrXKMI2bqQKmuOOtnwWt4+EuWBog7g5JEdPLWC3vg
pDIqn5sMP8Fit89JrdzvqKNWiVJp6nAl5+xyyU79C7Yw9Z3TLDM8CVx+HfZKubKT
cnVCAhxTZEEPThWo6/YHP8EzaePFtjcYpDyEAJBmgiX5lvmwY1B2y5qamyLqs8xa
wL5EsTYD2aebzMaFbYuzVI5yZm4i2aGSMo/8N8j0SxdCEng73PjcAQWxy39m66c8
g6N/ZZwK1CN2kWehjAjUfNjU7E1zVgAvlwXYIA8Sp66ij65vpB6fz7IP7ILj112Y
ryFEKCQhXe1Y9HjsYPgkj4zuPUDcyP73aZT5gmJHWZqxf1RvQZoM2PfiOOG9lDtL
O8Cmo+daDuy+SkFWOFO0o97ECoI3J1HBocIdO0H1ttxUb8iaGqjyc5iDYjh7eg0D
IPX3AbLobNHk6Y7L5HqlH1AY8WqRG2fptGLk/zoRB3rvGgfIIHcD2LSmQSFilQ52
AR+Xl3uTYMA/fh1GTAvpx70sNQkKXyG/yUOHMm2t2vsq0MJ1tCz3DHPc5FBX0HQF
YleK2DUGDPuMygb0cM0d2TPGCduOrIMt3vbrl4fpRTnbR+GlQziVm45csyTaNGcK
5caEnjEzhBD6MnFuks8ip7L3dg5Ib7xBi3zz1baBoFRBdITHEH2fnw4z/QXw+ttU
F/qsE1sGvYX27UW7ebsayK0HjlhSgwLJ9yNxJPyq+TkswWKnEczpBxmFlVfAv7w9
b6WHvV1e45/3FwW/HLrbztEkfC43xufkwSWcSIdb4uR95uW3NuXV7wTQm7fcBYd9
V05Y786N8zyB6I9xEpyEkxu55GLCUnaZ/jza5lnvHIqprAh3u3yg7HgC67tkaveo
GYaI8IRNheFdMRXcFbTuA3B9vhumhkhLCGOci0Qm5aGOppoTqAE5mzpzp9zseycQ
XaVJw3OZXMqum+aAcToIjIvqxLwatL9T1JP64BuReTf2ChNO/F4mTfDewo8cJaYl
KqKue/EZXWmCNodwk1f65pmSbXcZKpwMph5JPh1lc3Ri8Hy4kvZwuceyvlQ8CqW9
tU4WqBv9IDCK9dGHZoG6BVHYAerbG15QyiU2MhWuQ75q67yUvwor1xgkj3TE4W5V
hYnar3rOvE8hYXdut5uHNsZd/pAxIE3U/+0mlunWhHnJjUCwITS1Bq5R/2e/g2P2
DPeKyskKVEuBEnBgDaJrs0QbQj+k6iBsZn5UChiCN0MY3da6AZ7wsyukrlsJUl4h
b9+0CUHzylQIKiYny0RQdxf7hKUL+SPJn1TRxMFnoRR8sYMdazFQg1cfFejcztZw
QWZikzb9oPbaJRkiGF5oUiXVYTHi4qzryyt44Xji4XaB5lBLrIw70P1Lx6BtOTot
zvZzl4IM5SX3XD//v1zNaUV1R6hbcm7JqEUT516I8xUpc0/n0oEtGhDKLYG96Iov
drYIwSXlAdCOiS/pCxHRwQSfz2HqBEhomIvMM/YZiCdmcqO6Pgao7E1voMkHWSb6
IAiiKKZuEMM6gx72K6FkqvS96ntd6vP0osq4SyGAJeCSKFcnp1lLTzZ2pJ6CA9HZ
HCDYkmBup6JCX1Uc4RqI1zmqVQbUeQ+ykDzq/FvTpyQh7FhF3YoEjymMa5ALNffK
vOc4I/Kkx9Dpv8FVfVI3S9OUQs8V/nHlG8mrKoYP+R6wUngl2SdTeMD6JeSxlvLj
mVFCFO947H5bJq8BP9FlG1DIZPglmy1v5dMnDxWDrmxPEryh4PVeIAEF/W+wdL8o
xQxifU4BUomhLf/n+puKZtLSFef3I3zaJUxTFhQpc08kSxzP8KaDDmOJNsg2Wph3
2b89GLmFKFTesmqV2HrOyjBPWObbGkRloHN9C1BrwkWo1VB9T72oLOaZgFW0mmh8
1P8qsr7R9Q02BRaDPVR41ny3A8dh+4PNRfZc4nqW1/GEoFEA++75eSJ1Z2YaREEy
XqzcdKq2XME4GbATNHuD0LlXpER51T/O6wa14rvNLiK+qSCWgJDZTx+v4u2CaWdA
CZLZ0RBGiNj4BTeFnUb2QB22rFfP63Szh3cBG5KGO9fy6+psVknx4VsQ3pLO0811
9nRjdbweHkBrKQS0rlPBe0hr8lAU7D0UgTXzJjWbT9IKosoEHC/+ualBxNITTUn5
ipStr7IB0Bxtx5wKmxTY7Qg1nHs9aqqsCkzULkpX/kFbe+6DDlvssjYdy0adOs7r
NfO8xEY3GFZg8YbY4J8VWvqDOjaM1VzzUy65Z6R47+J0akpDmY/3ZOzUxOWBsMwW
zhu2GAO4dpofAMw1hlj8oJnqnJ214Ib1YO6fSN2Cir2YWd+LACZIv/bB0pbH6rWg
/RGmFQynTepqTdOti5QZWyD/YcAKjDiTA1q+TXQMr1bgo3Dm53C7b8f0t6s09k2k
e0Zyc7tW2jTfpgvleuSYEpzQ+Hjrx39/Gnd09VDuVCm6PBqr6r5kpGFjIDIQG9Sy
lNZltJloBjVFBgpjJdLEcqvuLAJZovAf7UcUO0bIDwzyRLtMfdlNpJbI54/Y/kfh
ooDwxdtZNyUU+419V0Y2YxI/aYRp905TYkxGAhjWCXj8rF+pMd0QdsWGlOsRd23k
1Oy1hkV8uISGdAnJY1Yw/8HtCBJkkhOUDXssPLQtNyWsv0vJ7nVjHx1hyzbckvxE
f7DAqtrMZAohW8DalFrdZTYYmXktwKMy2fMDJ2AKsUghkePBmJlkN/FCR+tcO6Sp
MhAV5cKXI9xTGy6F/KDa4J6hSPrC47nUBf+b0JtZ+sSf7ty2rp5aD1KY3DRYrGbC
2FtpjvUmsPQPItFaJfiNKyZoInrzymNN9dhiW4TuPmO4wr5VcmYsJKaOdjlwB85d
Qu+7OaOPxasBrxjVZAY3bIKYIxTidBHRJImuyIPTcO835/6P8WUY8SDiX3ugrqCi
a+d+VcAbT9nQN6IV8USlg7nNJ5feU3qpXzP58k0W/CNaQ6LrWC4lG0xKw23hlkcO
7DOu50fNMNgXbLdyaa35JMbwVW0Gk6aysMUKTmnD475sSevfbblhhvb3UXht9/R5
DK1OP8FhPEKsOzsivofxd0VctowzbRT298yE+wLUiZX1e50TFz+UH2eZkd1uJm/l
JWbeDk4cbeDyHSeezmt6YEgpKzsG2DNgiWE5AgRfE7YFH3eWgGplc75fcZ2Y4ayV
qzb1u5S7HdmWTWnwTYSUh4C7EQ1e2kJUhHvSchHszdTVqaw9S9V5TlCB99sKtEDQ
Yak1cMdIHAztnKj3eI2UxZ84aSsM4MUL/Ohl/YrImp8kC9ltZvxjjaeAL/ZfgBzg
NtJZ89IuwQjDNuqS3mvybSqnpk9t35C5iL9GDykngBz7zLySEElmuU5F707foERY
XDyoi85LuOXKdqfPP+GpUN+FCMBr1mHppn5CxrucHbjNZXaMrIwrEJ7j+QNsoS05
P4HkmXuGDb4hXnQNU7qJoovyCaM0PThh6Jqlu//o5lWrQfgJoeaFZeZ1bKmra++d
Twpce3Y/Ri8U0GB6oYPYZwdK6OAqTopcuuJxhngVbVemdzj7zVl2n8sNo0dHGnys
ZwAHRIZikipBDvaijPWmnF95kTaGWzaDoTL3za2jnAnzq5aIPw0Q3o7w4iOVVVsQ
Zfy5D2CCExKHoKW3q5eC7I1F+IT0a5EBz0ceS/a8RdlmgnVqlFSE+J0n+a9KovM4
O4vTrojqlRsMmhiFZx0nGTmYS4W2neEG7b+ljBBc/ojkRKQTwNmbzO67TXtru+X3
crscVxY/lB5p85EqCXPLht67yPrAbZBhUggSgHHUjYnUt52mF+7fTD9I+vMYbDfa
5i/vJYrUU62h3Jf2LxjJLsjPHvPgiVBFG4FXDL8J43Y7/TtKGWq3O+KXT0ky8wjh
c4zaoNf5hFRqN5ekCEwihBtOuOKublnxTijrZMJGfOpkZY71i8ouPZRThF7El4+L
UmRjZSas1tOG+jJh/X994EDCiXaSaCo6pg5o7wr/FM0B5t/OAu5qOAyIzVC+kW/8
gty8ar7T71jlJev75JjkcsFgm7hkM92ipW5RkX/JAnRTUqokV7N0UgfjuttpOK9P
eLRAt8fgJeFudtPCu6eUYACB2nTqgDMpzf/beE/6cwdsAKCG/aIWgOs8C6RfkFcZ
qjJit+9HVhjCzo7cCeakxTZsqmGAYxJBhg1UvOLjPPfGsRD9ScaTdZxdfp0+wnfJ
4/b11m5tBvvqnJI7qFCqQi4tydiQmsJrbC+ZbUmnXUW2IArZeqkuuohLn8PBG9M0
Ju0jxDxYxZe41s/UXDq6btE+uAHoJJmDzEdPUtDuvP8muXN3asC8iC0tp9OK5KAN
vXBxN6T/djzo5Ft3LrgN7F04dS2Ok+u2+Y3AScH1NVgfOpV3cYVjeOuyovPtg6Re
022UlMBvILSoSCrfnyPLlyzNTQ6wdVYmG4Kzwdf2c3DKNaZnzioaR03LPb3ozvNS
g3bsdXTsl1/s/KW/gFVPlvMa8hWIQoAUvG0/wLwaQPjR0KaVQoZMpBSseRxJvdLP
tMaHFoJg0mUW/QLA5AePKwYwF2DP1QmB9XkFOengObe7AkrtI5iNwIZR3grE/+bY
WN/HmO9qx3SJPWJysHv4+7++aDFJ5UWOaViz+W/w+Xxjv1qml/wNNqroDJzn73Rn
v9BMVXKubm2SA2TQn6X395c1mePtK+gyYte52uNKV4vxKAbuKScCE4xbic39kXr9
Zu2EvddgkeLu0T+EXktjgD2P3B/cvz08SitjOxiVfxrdev3nUr6jvkyfNFt9KUhg
b4kzP3+RMDJonxnWGXfcFLv2hruBomnz5oJF1+VVbZHjPkhwoHTtWvPBKMyYJmas
0og0t4/x4qiAMn0LGXQsiqyyMIEGK/G17bPM5CbUzYuThZh9ElHWgfUuDcUhrOMQ
m6vlJ4o1MLxsHfq2pVF8E2jAccBF7s7t3d3YZOt6XA5KVQwBrFj+PrMwV8ZVl8ba
0K0pnD8hL0wbex2SsyeSxyBW56JfkWARRTaT2/sI2nGaby8u0uSyauQhIuKk2TuD
XcQZ3CaOEbjCtyBbNAPOPzLml0Z49s43A+6PWEPPwYH0+DZTJAmFe3HHTHme8jHb
rT23CUUwj59kRafWZwifS4XigviVR5HVYTdlir6dgUUUS1zVss+/UR0GG1Xfh+MU
wlWv91Mimk44LuzIFuXO1JurAHDqnF2WZs7Inb+i+1cx3W0az/a4N7eqlH3Ra4In
s35DAtALYbQniJATFZVkEGW+U96Fl/LLy6O5gE5R7uvtsq70OrS9LFj7pD/6oX97
UV+hTQhSY+k+A+075QZj+SUOhBJvHFmTTlus4yFxeRq/RVcOm6enAk2+36U62rVs
xbOQsEEKR1HyBfEvOgc14YBr6qPnhqeQ2G5sta8L2bG0YFblT/5sqkZyI1JfRXtB
lRLLa8SfMiFwAQuk4jnlYQzX4Usz46MCPxZPDWZHI2lm2qJoPmSW7c9GwemaS81E
PuqTQqHsCD6EM1ap0pUjerO8FE0wTWisH1Eyjc1jfaioN/T+02hGFpXg86BZEMhK
TS00ByGZCnxYYFj2cz83Zt7p4FKRAfEJgUOGBDB/7h/kHHUFbO4EiFksF/MPAZaM
iosWuoI0kq1clRk1Pka42eAYr7WhOv6HJ+qUG7GN4/tWmsq6u6KbVQZIROcWGgw4
pxtbFfOmHC99LeHxlIvzJdsEdAObGVtJt1hbf9TUNveI2DtqYH0uBWK73Sz8sk8T
NAyAGTIndD3iCo1P7FriLlOME0jX4M4RIHznZ5VMvykUrUJvRZLN37JHBIjOIrvq
rG4AdQ+3iGWv3sT1iJjktR27jp93Fv3vWjzPoSLa2CLlShw1my9wlhm1NEel6SfP
eRKLXY+5bF7axq3EPa9n/3TkdFlDC4YTF5dEwyEWNSvcuWi4dNdEJONs742bYv/p
VDQIQp7VuRPAYVZFYCJQ+Pj0LhiES4EzDEaxuqSAsiodF+p19iyh1HV+ujyXYSdL
+phT8FUAkq8V4Zio01nVz0CzWdK38VDgO/PP3WgLbK5n0Sbk+jFRWlwWD9ioy9AG
m+1+o1cbmZXGOyDFw9DFvqCQL5k0BPIpi82N/BF7W3AuBQEy8IiAbJNMwXbZ8nzh
uks4j6HGkQbr3He2u5URb/Y53SIkOHjB8YBspNyCt5hZFZJzrxqAX9ZU8SLuM7qV
p9Si0yCoIN2sp4awRby6IL9vF0sbcBXXtDxoVCSsiViRyPm6z3J3UMPBmRyc88Dj
2vSrQsY0wujeIkHvqbTgz/NJUqifQCHL5sUjpxF9/EdzjYqcwN9mr8aY6kK1mNkm
wxJBfvC23lfvu5paov/+QZMJqgPJJ6S0Uw04+ffp0aktUzOx1iv8JuyTax8PEbgl
eYgxmqFA7LC6Dae5pnHYfWvGiE8+z4ZiGMae5eZEVFce1wwHVs+B3sgFmDCZXnm7
dPi8KMSMe32FjguMdDAcaHl+ekWkjfXRUPUJ0u/8nTUurxSWfjTYvwXnxGrlSA5o
MlGeZ4vTTIfWaH1ym+VLlJZFI5v/kUiTuI8FKMBITGIcAMmYH9enZEBaiAJTto6L
X1tBvyO/oNsrVTv/+fod6jYguRceBViBtt4TwjppELwWOf2vjKG8oqj18Hjo3aYx
Qy8sHHlXgvKX8RYaSQSX0NqFf567gJiWAiByzblZ1+rPoP3Mcxzb66JUvzlw6goE
D9ahJpULXmTBRsHoAZu1vSdnOTEw8QQjZJd0VbdSuV2DnJP1XKNVjDHDUKYJRkEy
AOfNl6p7A8WyF4QBckY2gF4zu050a9owRRb55Wle+kRTVUcGKck78x0qaYqPCcTP
K4Gb05QoCvdK3RJCxXVhGQRG/hkhHZuxLZHLTXSbH3rfQsNDb3kXnlsHuRiwswUv
rlNcxai8VCT0YpnJ6Lm2imX112WkjrC5DUnr+cZo/FVV3hlNgINRcaOCLtTdH7Nm
whFqQVSpnwzJ9oujH3c/RwFgm0Ngdnv8blGTTtquuIaLkIbK9KkqreoU8qLxtXck
v7D0uYZaJ7jyTGVBSSJ0F4jpon5wu3cpZfEVGiYcLUNMZtmCioNjDBiJ62QiYLx9
TLr4z5sbsPd3FdVVLstfMw45Km8fsIktk34DfwzLH26gwkId2yKCNoZ13+RG9668
5C3hpUXmdNGayV6EeRZT0lWH0wYiHx6Tkh/OgA0TpOhk1uBBe7/+GdSEnZNeYpno
CKWXOQpa8l0604IO3Gh7sQhuLp6yJ8Nm2v09u5lxHSozrVEGp4nrElpJMCbTtI7n
SxsZuNJJ+H+Ilmz3pAgAMhog7Ld1nvzLRaLeylYqRZeKwZvYOM3IfMYZlcI7ILAY
yRavnO/V/IA0JOEkED66F8hTtZCHW7onelLLS04neDDbZo4e6rhcNzJzr7X1yYQa
XEZ7nNFN9jAaFgWFwwuql+HJkbItjoq4gmWd0gA3+Ae/3cYSeEiC4S11EtWO85wy
xwo1UBinlpoT+5Fob21PALiax38qq+pckiP9zR0AMgvj/tuJt58aQPjs0fFxHLWp
KU9BLokJ35shwdebVeCYD2VLobZlYUm8FQYW9bFMlzgEFQgDHvu6iMUUX/96U8cX
hbffZjzTI4vJyhR9hT24zXwam0Sh5M5rv76UTyzsAPuO06pfkxJy8XvW3DTVct9U
KMl7BJdQiVZuuQcBFJiX6c4unDEN4efZjOLw10nneWu8wW4mwCXK/d835eeL2urZ
xd3jAFYG7/KqyshVyYwZq+DnG2ZndVDSaCmzVCeSkT7UumdnLRGlqKiy9KdBU14W
JntAcv6m3lFILjKIyUMteQRfxpM1n7jInd06dh9FZOe4KT9Je62pfZL+gWHU0ivt
fGwH72PPeHdBpC4IbG9dwmIipewVfdZdprjHNPddI8NNML2dHsUvjwsoicqs69RV
z7+CkkefVdiQ467ZJybMM181uZ6UDgiIn6TSKCK1JhDX4vZwUxsRPY4t18fYd1x/
+l+p7LXJZ1VuIifGG9QFMg6QzdiI3vbsyjwGNXefFL2NauAnlW0hcUx19CJDJ67p
MS/dfQkr0yQ7y9p2k5VbNc6xmRd0JGvgYrBm2OTav7mMiAsU1kL5Wsp/vj4Cg0YW
F7M0g09QPwEceEDjT7WZJ8dz6zVGJ6H6jI1bPotqvkbdsSNUtRPwv/KryyDlq2hd
RhCi7tlbKVMAfN/h9VNoUw0dF39+W8KXMd7F1irarGqY1ixIgeJ5xtOuYV8pFLF+
K1k5FPzhE5IFkXsspTSNqg7PrJGFaiKFu2eIPxKnDBkCwDTL6YdY+GTa+mStOIzu
TRGq258yZGkDflUUkhpwvED5aBGOX3iaY4jAqV+caRXwnlLte4uQglCIYvo6TrYY
DlIUtbY7Ew8Bj2SG1HIM3c2G/Sy6kaQqlapifMftdpEL+yfyA3i/C8rrVyjAFgL3
5BebTq4QvPVTajFJE6HzqUuTYWqFEmjNrt/nNJdZlyjJQg/koQb3IQUImtAyI+I1
dPXKahhDOXB5Grg9nHjw7wnNJZnl0xZeqHdJmpurx22DStwimJnkhL9wmPSPOyTf
HrpTGe8Me/mhPkXEVih+b2qnhFBKhIm5lhQZ+mNDMVG0PorRWJcrKwuXg3QOX/ik
V49h8KbqMpp6CLnak/8dELSJUbn+7L6QXsxQHKiX2UTGiv7fcBFW32mDGUlNNwBE
ve/I+hSwv8og8QgX7GrpcfbhGF277j5XWypNsCRQbm4mRzC47L7PQs71uphQ4vSq
7OKXQhcCIRX9u9p4pvbDM5/w/Kn4T5kmJm+Wpgznyr9g3maGpCnZ1uStQRu3jX93
U4+aJEjYJJaealMNh9+DnNaKBMz4LFCnMcfMoMrUXhASw6GXMMgWMpO64YlCBPYs
uucjUU0WrLljmKkhzDVY/2GqNw0g7wlinot4gWmRxFqxxC5XYXl0uAIgd0xB4qpy
d9ZFGoEEijZT0OkNffvT581Gv3ImiaXbvwEGcnq6L63T9Hu0oTrfh3cf+pC3lYPo
vA2vmI9VWiHUQkwOyRIkI4GQ0+Gb3j50vmtQn6ZVMv67qHVn9MPNv2FaNuCdl4fJ
xPlKa4JlDnv7W0tsO+Aqmo5hmABAxYfJsOSzAFwd8BvSnGu33UGs2vbLI2S8olhS
NeUxAFE1gx2Vt9qtNLHgUAhLaRjlcnhcgo6ZczIWTiRr9R83E9J/Fk0jO2J9UkGW
YH8IwVEF4C2Wofgnw21M0dPZhkHbUxoJAt6NIWbZOutxwvKih0BYuy53ZMcqBkFr
55i46Xba0xIDCRf6ITtsyXY9asr1ZO8CvT/hjYmST+nokMowQnfzWikNjirT4co1
nVLkir7S3Tt+V1DYQzSFpq9cQgRbadWgP2I68UvTywxtnjtGUO14gQ/NeEmx8gZ7
XnquUUAv7VFH6otAn7sPPckloi9M9PHWyHuj0ZkvEjodMTIqncdwSiYii3ErMv5j
gV+iIYUNf5SDp5qxw1fXhXfMdXXnNsrR8C90JlIVp/RGoBjbZ8Nx4Psi0iIRPb7f
olRuzarQgXxiEJx+sLq8qdZFLAczR/7wZR14WuI3GaRmMEMEURokKioTERkRupQ5
bt0vJqqgjApvtpWhU7M6ES9WRJpG357sx93qMUHBZkLyErDaP7G1hx9LCYTg9AzY
0mhyTbFz8Qxevo1kDZ5uy9PzEtnhVhyAPsr9KVwVBjrACg3CdV6Pbgg51mTd70Xz
VHySe6E6VAIyOcV8OXMpfs5hwmaZNfdYPJhISs5dFMdueUhwujQM72yb0QjPXaDf
IQBC3KdRWYOKNqgzV4t0r/ThS9i16ReokJM3uxbXap8mgpimZedHvw5DdvqQE2NQ
4zc+i+VtgQDguNs0iLQxgtR1d/ThuS6cyR+DT9j5vnGut25XWDoYGAlI6ggObdcb
xkAp/ZgPcINy0xKwiCwZGl/iJ/GbOtupe/zZocPR9Tfwm6UmO8b/v9daJAqTQAj5
brouifXLeXlgT/y03e8AYMO09lLpmAqvy9ku97BETnz7I58FgyehG/u4ngThqpqf
w+9J8mRXzKsDNc49ZJLD1UmZd3SWISPQXkpjP38aTAVHRfKumKClMOmF1ygI/2Nw
FAb5iCayjFylfd+IQCvK81WzguQWJQpPOn9D2aHwsg2TunL3SfVkeV/vLvyntY4p
b3vJH3V9DPI3wh/Fe9WpjTmzAXASoI+KXKzgzHZGi3UIw2cah4mNmvB3RE9Gku3D
HRgQ5s2ARN4+u3pwWdjCGHJk8N85JqdUvI32ckgSXtwhcMz2ncDm0pU2N0ZuA5dd
X5mv28EWyEHSG6DDoMxZJid5syUA1q6/loozg6DW31t5d139Tcb/x6Y1BujGBhtJ
gLcyboOaqP6E4nWpxdWVr+TNpZvAgEeitedDKGPz9xe7YmXgJ5Y6NtajR+fpSOg9
Ri9GDDOPKYWxoaDoqz0yQgTVQHc4cYHn5kdOXlHTnPKi3jBm1rFIlK8wR9tdgiqo
ZRAo/XRn1N6ovjy8ACWGxFxlanXRfD4r/fwhVnC/9BptLcHZsjjYvM9mIQFvkVbS
fdPNmXRZfybykjGO4MkJ3xyom0QGvchTcVCroQQ+rHN7PRBYUYZyoh5ITxvk1LOJ
WzAzkrRQk+p8mzIJawm1YYYKVYQ7+HA2QLt5YL/hBNHhHTpa1sZ6s3xhz6H0HbCs
gbqyoLuwxoY0JzVde+2Eid3Bler0st7F8p9ghF7EEhsr0B6MLQPoWpeWuoypI7xj
q/jR0SXWYsrNo30AenHDS1zIOa7kmhymeWfnUBlRaKBCOEZi8XGb0EmT8jnIK94y
VDunUmk6GGDg3mtyYk8UdfHWK8xRhf1dR00G9IwoeXEv8mmYuEemC5b+D13OxJAV
/nRKREovruXxKFTAjaCOrKkjmdUevkQh+OAZQcFCAGmG1iA0SvIoGi2mnR4bybt5
1phTOPcLNx2DKH6em0pzFtkjJ4VmxEQfYkREjOfx9yUxsnPRUDSyrLfaZYdMXxey
FKwuMKYGlcz1HLGKSN0G34vwIPhdZ2bMZv1H+KgwLGyeAUReSpp6/xnO0GensCEb
85yd8X3JBKsBOqV71/9yD1uDFZtemb4AfQIIe8oa/wLpPKEUB3/lQnNoIWA/PF/A
raAErKTZB6qAG0TAIywhhqeKz8cTGn3HmAi5qorWe5cWyonouxCqsrjakN0n1sQq
BqyekUEprKznfYZsFcwjAHzOtU0Uz5uyBAehZUVpDB7tFdMco7GCGVUgwV3psebc
B6ys+BLy0WWhY8lut0VA7c/hK7uq4ysUt2zI0WfPCoOgzfklPO54rOvMbSmXb/+7
5Lg9hrWxKkz4yPRP3aIH27CIRR+NcdD1s7tnF7F+qQAfgvYz34leVCG6riZ4SdEE
cKXF5GtQOUYjuIauzwu8RckEV0Woqp7zfsHmyZk0CWIwAAi6xF+Xo8st2GHUFRhB
qX3Jke3HPtdsyMh8JEk/Sa1FTy014aloIiKO4/UbqO3apkfiQRPNTcHyUw3mggAn
wcPHXogE3AFjguA+yYxAuoHD3l2TIL1YWrkqWtRWnk3YLI+hfl3188JloTO2MpM7
kKuRX1eI5gYcBVHEUb00OCVrtX2SPdDKKU+PXyB435B6FoQLgQer+AsmiQJxuVeG
GxYufC2ZcU92Z4KVOMpRQBPXPVQk/zTmp1wI+XrvU5BMgt2G1493Q6shnVMOCMXx
tXt/eHIP/Rec8XPOA2P5zDjPCdAJypwL7cB2B1Z/MxHIpC4SnAH+9vhC2Csecci8
xBw1p2I9vbVzXe6JDW2kUdw6ZY1fEZC+oftdl4i+2LM+r2tai821EucAh9G/dpbb
3joXTrsy0BRh4agvfDZbFVRlT1B6ozGdN6uh5dsGSIOIZaU4O4ZRT9aHXYkohhme
5mxiEuKB7sGSQjNbSjhR9BfzIDhs0dIf6wkX++IuuGttbPTIAGwNx2MAHiycR46A
C2XCsC2mvTvZfqYjLbJHK7uuUQdozAhg4rFGSenUJa76g+cfPaINg3lT2c+PLJIP
djl9Qo77tWQSAGgaIrzAC3079QSuS1UX4VxmsWqP5heJjneNOTSZEMuTmOKzrZjd
REYjtq7ZAJRS07DyfKobLcj6Pkm/et3DNOwwaCIoe7CGOkMTagsFDun2DBtF1EH2
SQbd2QuTnXokwo8l6ISeCe3xVGMp+QtRIltVcRAdBjBrH11Lped9eJFlsq93Lbgy
sRHRN1QTpmHxpbEoBT3WrfJ3PlRdQwWYDQ9Io3R4d5ENKsF+5lI+ktTVa5XEXBHf
fA1SkQn7KSJPC1c85laNVFfzkCFBtDCKuhIQpcyrigg9mq2KWQgMBc4/s0+0xXwN
zlXFFf+xlPHRb+qKuynUsM9FV8KRBuzaVT51Pwcnc64SkRc31A7H+pcR+cvw2Lwt
odYByVt9wi7d13gNfWXVjmAVESsEii/oAls/04WMOFoSM7J4rA7Dq9Cm213YhZ3k
a9BThFobsnSh9rthfKLPr1oDktk87OmQa6Z3z59mbMLmKk8jOEUbyyLkhMG4Iafx
oM8Wn4VRDY5uNDPKkk+c9JljDY3hwE9se0bTUSyeVzVDpOLGxVLWR2U4iGE/hdjb
TxFgYyfahs5CQNY5/xTiuldRjCP2/ZpFXU5ZabJIOXmq7ZlRqTublpyYZfMt9IaI
99ZNfK97eHDGSWBOfMB1fIX6ps8gVLodrhnCHXNan0ye4KKfe0IEXzHvnkx8GaSF
2mjkhxkXUv2WzWHapfB+awmiCaKmX45glYTOSzYU+9P884Q9tAfc9YmYY5AHxLYk
fj5TLoNYwcByhlO1a50JKQA3HBzubdcxLEyYWI/+iaZ0YM4B1ONc33IG3EDcmA34
fOoZ2/osc5oFHmufHS+GadwZGCnpQucXPN8OpEVAWd+aH07Wyz1yil4/Uwy92mBP
H9IUKj88QIZQlUDx0yRti19XQ+x7pstink8i4E0oWxdokU7Iu2BEGIvOmi9ruvR8
HAfR2C26JGEV9MSH67rKRG2jBW4tnON1TmcXp5UfcuSjPf8+LY9aMM0YfoAtV2ZO
etqLE1DMXxR9NtwNPmG5CaUPRANUppUkcmqQ1y9lBghuL1hLJ0t1pV0ey/tF2PfO
RVRXtfNmJAUtdVCaaLPYpZG+ZuS2NxZ3BysvERtVCYM34CXWbe9OkUpT/xic5+Nr
iB6SYv4ew2GtmOVwZCot2gs0xm5VWCnGLBmvx1D+dGDapM7A1xfcbvNGp5wsHpHi
16kTjVoqEajakx55EF3VNqopORnhKk9t708StU0vL5uWZwBpNRrEsHLzwGQ78K54
Adjw/h8bkXgzABFrLda02coVf3FPlesrR2TGeh9AuAI5i+UBy3GDAHTbb2uQNCWJ
qy7Koo3t5v4hhIMJsnxmiba34xECf93sQC4po8eUnKW9R/YgV9Cbis6+KcEqQe1b
+yokiwtljYdf4Y0MKbtwCcEU6QuEMWdXeqb4LpF2Ldq0iFz+6FtMiS9nwbXFAYKN
YFF3qoAkOVocuHEF3alGIoOD3VPNNUmOR9VFPQSLxjML6fjilSPfOUrYDdjjrtJN
gAJtPXPfvKcsADjvasUKLFznEBVs1vlMw8lYYJr+OsCLYwyBexIEBk4TLU69AHld
mglUhRyaMdWsbVOeLOj9zF4jD+KQvVYhiesOTRPSS6cNrNPt350qqZruGC7CUmUx
Gs6IQyaPHFT7x0P7qaq5rLdzf6VsaSyEWLSJGKmkHxEXo0CMx+QXZpYO7z14d6hQ
ejxsykPPFxJE2wREhvicP2XMPizPgMUlJ/WVN5KBPxl8RaM+bpDuTW63IrAt4ZVx
JO/v9hGc8KH9/dghCa+NjMas55TI1qbFZpa1LdNZtQqOddK2LysOZSyDzwJl9wy1
bAhcKmRVWzcmG4ED1PtWPbM9/NBOWHjhv7Q7wsh6rbNahPUGhTFz2oKiCX0USxNI
idtVgWkgwMx8GDCW2FSG/33OS2xN+Bli9tYCirQTKzytkPphLOmsQaC+/sKlgQJh
lwNNsTuPW4mv4jKSoks/9T1rxYA0bIPESVo6yYqfI+MQAvcL5txL5iVQTjZmKIZN
L6fEhIX1/Ru2hHCYnCHi5O6j84bShYjy5iUXNQ0xRO9FyT2tmkSxRue6xEKjmdxr
ndMuYFwT0LrGVwNTQcs9tU+dycStHZYcdb6heQjT49jDu4CXheDGZ+/2PwXZHi5D
6X1ZpeFyRlGcgu8lBFC+DQAnUZ/GLa6xaz8Qq6LVv1FzkDb3RhuIL+5TLNfQJ/Lb
pVpzbBPu7zf8t4t/ffKoCZTcPhio/3vpbkaWatk9dVuKYKKm1ZfFgb3/EkCYDc1J
DS0dYWbOIYNx9x4wOB12KEWsmCjKPwJm61HSAybec6oi28ymmRReTtk1Gl4xIVfa
xm7tUCdzgf4s3GyIxGLdGIa7ChVP6lj3n5MuEFpgCy3TQznpalJT3yclJ9dUXwK3
QA72V1OrYwQwnPw5mO79GPrxCJFU7Sdvo/1YMV5JuQIlgyKqhv04FmMwC2L0yIbG
kyAMj4ICkwRyYl7uAI+Yngc7iwtcrm4pljMaGWm7aACU5OFG67XRQkQ9DetU6SbN
m7PViirrIPhfHKa3+5Z5pbUlIHpDtnHZ+jAQtSZGiD1K9zh0sN125tMNXNJ+CxkO
9j9z5psqXUzi/lh3Wa4uGA4Dx1DelUJcMi22QYkneciaATc452SZmBDGAIjjfDYF
jwBRG8FHPVrzGHNpkPSwF4sosDKhvkzal0w9UUxxCi1crbBPW76jKSNqWGGkIPkM
RomdMFd7WG0rHoTfYfog/pknS8Rzzk4oCb9OC5fRNjR5J+bnUlfbZhYWfbbVRaiH
Oh3R6foM7oF4Fj5ysch1oijHtubk5stC9fb62OcIKdj3SNQESGQua4ww0Ag/b2Db
31TxhxAax4O3ZQWu8gGFJm0L6E526X33jsYhUyy20G3Q0JhfprWNWB0Z7g/0ScKO
NfTTWd3V4WPBjWHfIX+ixyh4u8A6hew5Lp3c8jOm3Yxk3tLWhESjn3ofdaSpHa17
IsYBgAYLVB6k1ZyjhTMa5x9+3wKcTVTg69EJDStH37ScGPcpyIeKh3TujNzPzWBy
Wzk+6ES0wC9ArOAshPhQ1IOE/Ct91b+FY0mGDbea3dXPS32VsS+chlptBxL9ZE4M
LjdTxTM9y22FaEodStYQODpj1Ob8JBhrcUb6HkqkM8HF38y78yWmUJd+Bs7jd9cP
jWgObVWMA3gKc6wTryyvudq++cE4MzSIANbT3DU2kIMZHCEkluMY0NKmnwdj6nLu
Wwf7/DG/RzrCR5RhHDFHMtRqu0RB3lpV/qsnH0bpOr2C0xjAwWiJHMCwksm3hNTr
ReN8my8A9lA9oMvXKpdkCKF20aMTd0JBblUqvAWdp5BjnuBYUk5DsphZkdjzMb4x
sUgUt0qlO3mioors3DrDukM30yBwMQbDcM73pMv70xpB3erRb9x1ouQqnYOeSUkd
gibcHdsEC55Pb6c/OIEMmd9z1eySFf1xf2e9nNL3KlVvHDnmJ5m63Pfjo6KTCKkB
Zgtw5p46781Nsu9p6DYSOCu2jzcQ+qJq9Ybs1L3VdFs0uNP1dwjuda2ajWHTV4V3
qsPsAfCHd1MwmrneBNfqz0BuZQQrPpE025MquLUtup+9Q0i4PKHQZ6xfZZk8XVwL
CbviTihov53spjfQ/TizrTIvjkwoB2i3BqKiuJLeJeZJkE8zyXugY0LSYUZPHfKf
DcjrQIdTit8ggpaGtXT2kh8qed64DSAwKZMvh8NcWQH7qZZysakaqGNEskh/dXqY
uVzUIYrvRyyr/KnhIiLDvHndDOJ67iStWgG13dqwF73RjsxbojUVwnv9bOoGCuiU
dAm4K6yLIeZ34/1njq+RqVGyA+HynyZX8l4DJzxsjGcPfbJEuONvzIi4bFOSmvRR
uXt0kqOCW9ps98UmOi6Y/s1tuvpvc4gpRNOLI7GVl5rGhAmc8w1zybq1fuSfFf5I
fsUGBDdOP6KK4UEx/+46Ruk7hsd696TvMRdTggoetYMC1iYwrBOuVYlYP7oWnTsT
QKto9I2uY8yEPWFZeunbwyV8ubEZSkctR7DWlO8S52gXpV1VNQVbDYDpBMGCiEN9
hWIDB2suJTfXTUF2U3qucu+KkDnjaX+oGFd1BdgESV2R1i+dt4gCTSxEV/ofxTJr
urneDO213xdp6ip658DblW8oB7fyzmb5OsiQ/Jm8DoEHnDYBipQ4RLpmb1q2NciZ
ysUuNt59lNa1KZumVCBVNLz3PISik2zpHoJNOVsB7NFc7LqG4v9yxJZYLmLXeefc
gcYDq0m4uvyFwYtWBnu225h26z2ErDdDeuTElKtA7t2nPYvLww2hS9fU4ybs80AE
+xKeH7OysdvxBHIQ9vftszfKkkArBI4pWatI6CKlM4ow7yBwcwPFRqI7w9D5+xpt
SLtkdkwkM7x+LdhI+j3SZptuEtSfHsWBTXBNFJxAq/UTShN0h4HXOO1VrUaY6Gup
K5e9BPjvQyIHJ50NrYToUzv1ggtiUuoZ6aOObIv+AKOPBvVlxM3ew3kVi+jaVK6a
stX33YF+ARUfWTnX3yEkNByKiDzG5r0Cl6xz1x6/G51OJAQ2pa/Q/idLUQBLmIjx
21/hZjmRNvgR2Xxsrm6TrGYV5bHh/6NcvxOhY6GLXJj0r0zEYtvOCvkfC9wTvjN1
0tJ6Ga+oJo4iWAfdJy9gi4xZjDufD277TX9wcq/Pnd0gNECkcyHLlkrGWoPty5L4
GmRwJh6iA/OD3uz465/nXYQBNhguVmrOY1J9U+C5ZTzxh0LqchwAM1NXaVdDo1OK
jNeZEuIRrbWV+bNzRSIGplac7+hjMGZ4H7Yk8L8NZcZz53obLZ9bAoGtM48Lan21
VRCh1lVgGBp+PAwpQRPPianBQRUs/TEFZZkg6QNLyZYadoXWHMZu30lQ+B2CgqaA
qTjYtn/gAd/lbcX4PdY6Q5/S/lW0jhh6bcQeutSdN3mcsVDwdbCGr0//BQklfWPe
gGwhgABuAgVzsBkjoYV101RUKeTT+9k9NTxyo9dcQOooeWS/1VgysivwpHt/phSi
FFATPZJd4yqP5VDfm77+f7vwyyBoyWccm/M/KGHV7jxGYoGQD5pE24VuzL8HezvB
6eITTu9X8H19piSo/xGD8WkU6xylm8YkJpDAmjs1k8K4KdEgvloLa36PzkK8d87v
RUVcJw11tLrdRYHk8fdwsTBUjK7DJzsR1roo0Sta6+1e7DWvd8WVjRh5CPsSadNK
MhCg/eczMSYTytmd7SYGuZk/egAA04Z8jPEXcDkFed+EO7Tbw1oQvmYMQ7r7W79l
g8dfL8JaQ5EcPlkJpAMHT5LAfPcfdv3ibQgIKkayez28+XG+qSRrce4X8GEPJPSf
LloFu6miPKxPTKea+TJNwh2vpUkRsBuOtKQSv5D22M7ADoOCdIaJTdLJKTcRmrG5
QPxqGaPLAbo2siFvqIV0ZPjsQkrZZIMvRJfx6UV1N5YwBmdqSIVHvtE/sxuyXlj+
JXvCqsKhLPfxzEFaxAosj92C/wT2+ZPqPWWEpKk+nP8goKTbLNyoSh0OVbIvdbqR
S8fUR7HU24gekQHb3rLlY7ylpGAYbrgM72igrEjR3txeIN3HbLYXE6eWf+/mayyq
74YGw/ONJ/ArjxDkrUIeTG2jQj/HjyL7OTqo2CkInAyd9rqNQh7AMtMyzk9Kj0LD
1zgg7kv/e5HlXUErkOCAa8Ye/to3h5uFL3J0DPhve906/ERdBglUlBOho/sCL1in
sAZCDlS2SUE/qekgJDUKsXfpksssSi7MCap5gFiNiUXcHJxH7uZPVuFLiuxIH42E
SWmbBvSslo8BxBkwGURPEa/zoJC4mXs3Et6usOQkIWCgyOfGMgd1uLd+geATPnS8
1JNxIGqqPtRwTL1UEAJgCaHW2zTfuMnZeGVu4rM3olLCJPFVGUYyG7ywsCeLwWSa
UOXmacWvq/bVxfbIG7UpAHK/kMIlH8eWXDarrGER2u45Goo6CNuFuXfwW/0w5FTy
nwpC0+E32QtNcrYu8c1f1S5n08OS333i6g0WOeEVCgUl8qY9su1WJhJ46U2RESUm
02agC5kVESMlCQD83yBWtFddrGwYGbBQT1snisTtJ/p9/ntSWIBinjg/Buc4g5Ul
oWEscnkVegzvx04oFQAI1obJN45ditxz8x97HeH3os5DjGE+9ij9KMY9ViairdlV
QK12Y1Xk3V8p/s10BMaEch2ShLlFXKX6LwqYC6CkxntbPpr5wkVGOXVu7NY6lZP2
WXSiSiZktGIizUiYu4DYXuZrm/Pp5q33NvqnN0AXK9r4Lj6uL2KOMNEdziSdcY40
1N2oChn3Ayo5Yo3zG1wm8LruhYG/UXIow4FTgc22L7Wx3EvYcXnc2cDCpzQGy1pb
Kg9jhkPIScDLnFPNlrqjDFflq31QcJFMaoWHOSiBEReqD8vSfxcm0cNwF8zq86Qt
osrS0nDBIv6m+5kMKy2h1IqkFIV5g8lvir+cdKRj1P17WyAytrvx+696usHRBC/9
FPQbrz12Pr1ZY2kU7eNuCAHkBJUKUhUpgayhwFdv9r6FmmINRS8umrfNGQ4XCWcP
JWliV82I5VBk/00CB9pqZ862sn57pJsi9Mpa/9fUl03OIC9rcXPvRomt+TAW7og2
HxjAPWSVxIQ+p7ULBeM3p4OAt/S8i8DQb0oObmXP2lAwGBm2GCj8F4y5Fv/bRWeu
EWZkxwZ/ahmmxLXQ8tR8fgQjDAJ6ctudUOMXU2M8Iap+4Ox/oV7l66F7lKZhACNk
W+IaBPK6Q4lSAJdFbGCj2X2fwDVpPbDrgcVVKREB8IIYC5gEE2O7sl8JoaA+sAbW
YH05XniMAMoFe8UZVm1lmPHLJxIhNgBP1sbbq1M8fMvpUUigommMv77ifgyDYOPp
Lmx9kMGuKu2C5YNW5gjBbt7w14tdmWUeHzLSkH4EE9iIK7NQgxFHeoOhP0KD0h3+
hei2bKxBiDxQwEPVD8c+70m9/+BANRTsNuYEBaTgcfMp+w3QFzWf4ghJhUFNnT1Z
QnQoV3J3GAGuLb+3StQZ8fPlyYhG77+tATra2nWUjJjp0nuLAWcsKn7yCkSh5KJ1
fdbECqeRU4gngpttjoglHOQhb9FbxImOJSvk03bC95ZclvjezJwGTosPTjhOhe+O
MWvPADKAhynt2cw31T6HdUuvEY0UiPJk3YCt44m4ZHSKTun4X05GzaHbnkMAJVNy
KI7YCj1vFufD7887S5TvX3uRet8bzT6Di1P+OJWVNHoqYNNx7ai3USP/L9uEUU5E
Qqcb6ACUqwRXovltCd9akMTxliheRZ9HioR2KtsQ5Gq3QG8ZWRwjDytI87mcB765
HvjZTiXe4s8H47EJqbEm7i/FPkrsgpRPt7F5CFk4CX7DNEjYUHI9YywvyKrxYkZk
MC6ET5OpijusKNRhhUO8OkOuD6ZsmIZf1zY6i9+1KxC7yOmSY8iKnbH0Ql+7ctCE
x/prUSb2p2B6IT0Yb1iW2cqGo9vr/TdOx51uxLrFEYalXeJ6bnGNPJRhauGJejXX
n/339UOb1U2EVCz7+EnKpjY+dLEl4fr4sAxMZlnr3saFnC3FMCMD24GFXb7pB67/
zc33BOlCNbmg2N79uhMVV1Yj7zEgbsW4Yuv+nZEr8sey/HvyQL/oh/PXLn12QaZC
Q4xek7vNw4XBxjc/KYgZljubkx+vkWeQ2AD9gdTKVr6yRXBHXwbMOJEb2K3l61DL
F2TE6M7MR7+prDB3ln3z4nPv+n8AeJHCYdD6lPT9FxIRSuxuRntzHg7dKp+zit2w
1ObSZGEaMemD5yuJES+k6hCenFLT00vGkNgDveSTafopXtT4frtyjSqqiHtRNzcL
LV9fVcQLn18QPVMnCEl72c9X1VSt82HpKZqBNGKwJOML+u7CR6TS35iSX3Z6ALk0
ttNjIkBS4pDQZrmNFTRqxgJRwnbMjVmU1LBylPCQqTi0ioQ+ZFfYLjk8uoIHwXcq
ONtXDlpib63aGQVl1QNkMBYxZOb46Z4q7DjEEmJR2E3PoUEZSqCOnL7k/CPRQidG
LzR9K0u3tiEiCxyQ9VujdHecxw25Hvpxq+bz0oe8CZF2CA+HRdr67ZkzzmAwTOpa
1exU+zBDAPbACTljtjhiG7KSR2nSnJN7EiVshw324r3hbHMFa3OJsqq0cHtMrXki
GsqJKhqGxGzGJkjSK5kxxYpQkwUWAb5PG8VA89JNW60spzeUBtJVVm5iptV6KjQn
vrUaOGBqbeKEoWVEWqXjJQGAtgU7Q0Y5Z5N8tmeKs/mO/dogsbPW6/dkQBRqryLk
YzYHDqV6O22yl1u7iZCBJ8eQ4czdRoqGspu1Ls5oz+/ZH/VVYJMpxlSVYiunLDcU
pBlWa1rJXhE+y9wV1sTTO2pBEFR9MF45nkDe/X2hZdQNC/OMWWiwA+oaH/v7rQB4
dKbN0Aaie9HzWYJQC6dt5tjPTpSppra1cM8nG6g5M+5sJzth5QPUj5mPiv8G52XC
5H8pBYTh1ztPY7UX/BIP+1GGPoaUgSzESNa/olINboIM1vusReCy5nc2RKcv/VIN
lipffHf7cjzxk85WqqzYxqIW1UQRmySl2bO6d8FEKxMbQGUY4hH06+ttD2stxH6f
I52lTGY7wBEvgSYEQGFEgMajYrViNf+60/BZwHn92vsZJPbbGkS4l31+H6vCZj3E
h+BOFOkFgmiaMD9/+XJP8Ay4sKOLpvcgrxE0WsImmcLurHaMAIP6UhuM90oaAnqs
2wZ7vz4Is3ZKQdbrB8YKsJS0REdsVl3Nl5ohOJ2729SIGECW7B99ve36ZTbB3GPC
+LsK7UjuQ1TvPXezt1yyVPRBqqeIlCKVVv4NDZ5RnvwT0qMd+9z33zyjjtwMgZzx
8VWh4TtrRc5FO/97D+HqkY+aPWk5q1yQhBDYlBmt9HWXxavwV2D0c2/5HqN458cv
RuTyczMaE2g5CKaCtOoGsagTS/RfI+5qxuztN51t2vKKzCNMP2tOLswfNLBdVArc
ayBPd4M9coJc6MdOLBk0asawPoqBU0Z1fH+OMMh2FdKRT27LPW23qm0jB2eO1+Xb
n6xCDbZVf/O5Phz5xS+fubYUFfAChVdw9HvMH6qufSv81jDx/LJ0h+AlICQA6Pon
ptT2vks26FS6QM+gAnP2opR2Zc7TVKzRelU+XExP0l7N4B/uw61Yjh7neHR63WIe
VmJbSv0cvqeAkUjJMFoFavwfs7j2IHZSjRq1LkLMhIBuU7z7v66Hlp+oa8C7OAil
mcEoX8wItqJn/cKhs8X0vhnhqaRui4wx4rkCFC9yrBOR93366n6CLHBLYoSZoB1L
/NTL5LkW480XUrGN6E0jrPAKmbq7Yj3um/pwebBzu6aipy/VQU8g6r+pg9zT21nv
ofq6QqfOKV0bHpYsC0JH8EC019uZntTr9EabQOb5AzJkc8ZLosJgR9HC8fpSQw9A
O4Zto0OaeOA4GDAyzgfPgq0cjYfpn4d44ryaZC/R0HS2V2f30D0Dpnp84PfnB2f4
ZWuLVMz9t/dE/LM230db9tDcC03DXolBxz0ewSenr8rQ/iBlUEwWM+kQ2wpZC4wk
nRRiaOrJKc70vHiqUYIYrMpfeRiIHDtLpa8NaDZznhL+gZ4EtCQZLena7FThszZ6
duqVbs+l9TuMp76pI/C85vOmZ4qEsoxH7AZJV82S7u5VwnlxS6TnVNE4+oVq3JN/
a2HrnYgSzS2doB1mVCJgrk7oWq4u0smn7cB6Ms3HIVqPJftR5bqfzfa9Tj4Ymz/X
5I/cG4aCIbB5H1tnSuiAEQyYVH2Cjq6bI/sO819rMWkjVxWD+J/2frjTI6u+SEUk
DasBvloSjhykye0705c11n3tzF4TdG1RybmsYql1g8OxjV13dxEmMXjHfEwAs0xg
3OfIt+irA7z+Y33khbwmShYlUMFxhbuHqSpZ4bCduuCecQ+sAZ3c0Y2LVPVIPaAN
d6BHPJ6AuHYR/2LJGXnXEGDsd/Atazj3Ch5oXzc2F65oZ0LISy6WtzD+FHzNb/98
mQK+lkHCGWVS6+SFIxXXk4fDsvBUQObveqdy/9FhLoaU7usTOSjxlA8OX5a+4QfR
nzfgF7XpcsmF/iI1Ka1QPRRcU/RtpamFyM0sTOy2ORCD3pM+WLURpQQO5Bag+or/
0u2MkTbkaaNWGHAuUFTiqhTqWQdJKGKjvEAEOlq4GUmJ80VWI9a6o7qGK3IoBpy4
g+njXt1H/tNTBb0VxPRyeAA0tfSlsCeVp5U//2DvN68RSnMQl4NkentXY7dhlC2O
N2P2FKBv53V9D3RndMoUNevrmfEU4DS1EBl+gEUM4Ed8QBOy402N6sdv58eGX5PD
YkJLvs6YU6sBacr/3R7ttsqA6wZ8Xd9F5GDcpIhck+ueS1NpB1BCQkLEybhfRotO
4mk7wcW2WMPVwXRD9UHy8BkRjmfpg+/nbVYDFEJ1uu2GbL68jbwrZGhv5vuYIBTm
Jtd1Ow60CZIJVKByrFDOHcunPjYzAVDR+uyq9gaFFszqjQUEu4ZPdu3rfEb6AUXI
tZG4NLkYlebT1mjanYEycPYPbki3sgg2qSVpH4nrVp90y6RXn/Ef9aQY5Zkt3jbN
0vgzVGQnh4LTqT7XiiOBmTtZsx6T8lVJ8JLnc5BOH9+ewffLdqGhBR0b4kLYHOoe
zkSOvUZy/KAEMoBvSv7wNYB/MY/FlFicMs75NKRChwu7IqH+XzpfsqUiAIjtNqIu
R14JLiKCf+MyXL7EUDatE6KOf4yoJ4uDepo62CTqAJSKBwJaSI5YbElJ3ix1gXes
4goCGC8wr/rhVm7OkYZ6ACQGWzCSlgAUNmYNwpYwN01anfaJd6Nd+YKvPZ+6rFe1
kGLQwxSp7wdET1bIYGXEtfKfqgYdp6x7IleLF/ivLw39+vDbhAFxoez1GJQqy/nO
8LmHH3TnrovjwOlvGGmBo7AluHTXx/Xq2jCkDo2pSYYA4XjTbksd3uaLxsJNeGpk
0LTkYbEewUlyqiG7GEaIVrhCCMNn0le3vOjAjLtwW5iQXNvxUcVhVS5ejFqvfrFR
EQfA3W28wP6X1VEs6QNhl+memOrdU0bz8eGHABXX/awOQdSyP4f66+FyTayTbdcy
e2b4DeNzABrwlA9wYt+93zYoWXGP0WsccJfBpDq7TafF7QEJ+ad/UKDqrDTNKLS5
HI8vaR0BQ4A6XaD5A5FiRSwtEgWodr5YIq4YeGCrKY19CnUAHC3z3q4EGvo3PpW+
xdfwZvwK2dtRh7kEuhXprncldqYDr6kmzlNXWPEscLCXKC5Q9ajlcJcU4Fy54pxq
X03bB81qv8PMDZhLFje4TYmgAXWfxzV/gNrPf0VJpzPC+UyqzU+tgrYk2i21zez0
Ao8VDRZdhchY71ABwWFpCjlNIKs2VZGUn72x6I0NBNF4fZHY9IjVqivPf/30AR4m
4BVqczdngCmg/4bBsCnTngB6ULuPOFCCirDHLENumkZndwgAk2PR3lIjR81ApLHc
y8rui+Xbf4cJckjYC2+dC1xjeKwFBImzSfUGvLTa627kdT2EVYKBLlcefFFlbFI5
OWLa7Y5tnJZk1TIYmwXVYRaGDGAKZPAk3ng2bENrF//QK4om2loqKM5OyhFHapit
c6xazN/vI1Wav/22rqM9Qf235+nYzeAMWN9U3mwBUhqw87SvdYqhRqI6XbqVXmhU
cPOtsUL1DGkwHHJgDTNz53FL67UbV1k8edh/QraiQPVVdrkFPXSIqLetJljFcPMQ
HE4kkqc/DxlAVjh2Q+XjTc3W0svOrMX5pAPHVLJKZMv+HAnIFvUMk/m0FtrXj3hx
X2rGlOCzu6nPfw8Sc+jABj/TXdPMwnfHMzNtYon9bMv9FreksqgeH+JqGwtRJH2X
CHECZ/4a7WltODTP+Eyab6b4a9/M7WiRcBFawfc3JKQz8khOmjqt/lTrqa9q9HAm
SWZc7VzE95ZUe1Qn8ifKotk1+FtXFzHCte6kp90yWMTdR3gevMlO4HwhkfB6vpSd
4aTPAoq5YdAo9hG6FxN2gM2C0qMhfj0ERD3NW1oYRGXEW7BxFLQT7L04yqeG4Ytb
IQeXWKZPVPRlHP0f/DGrA1426RIVshNZzJjqHoRriQrczE986EFfDvAT44qIr8Pk
In7JFjhKSVQODCEdTWCxu67JCih4Y7aBloQ4xaL+L/NVdViz93ewcuAhQzD00Aov
m0XhlfmDq8Fdl+QejDzOucYrKYGFWwHLXCiXMabyjCwkJ6XttIzX3k8gStvXpT/P
JFR4K8sSUCm/UaebWGm/wtxM6u3UD13gnkiEgpmZ9B1eKI8FibNH+J8rAZ4wWUW3
3ykNlRs5+0GBoM0IBGtdwQbbPuTZ6mONRPXyT3LI0Aet5WwAJ8jke/yBuFxkm78Y
ulyQ0igb6LkgD/pS7Sowf7WcDYxLEqdWXKYVAMLG2UYprvSuADNl3oNr5maH2nbJ
qOmKROXHixItWBS1hFPYKEKjpM4/o+R74WWB0bghBuS/6KxEXfUcsb4BA+7fB/9w
GThgOhTt7OveeUFZaJfCeH9fmncdsbSoaKaN9QfAYQ/UbBNllCMDUAlwyCAOYZov
61H6qwbHCp7nOQIIDgVJ2ltsLGpylfw89QZvgw5BR7yF17xyoSkJCUrXalZXX8Yh
takeUHb45SyFdusu9w+ZSshm+uQNmCX74GpgOcXNlIMNXdqLXyH3Qr9uuViTzkfV
au2NsO/r5NlGnqsoJYEwD3cRr0XMaoN2N7/TKemRAY3Srd8I8K2wmBKoi844RqUX
F9TKCA0p9lklxRfjhbthk/E6O9mvJtA3Asfv3NVuDhZqiTtVg+f2LJRNMZWhjQhN
EoO6vCunDl7ZFB5H4qjqqeK3dvVSn9dc/HvlyqoGEsMq2pS7FNhE8ZO+LLP7DKJh
bPMcipeokG1ttcuyY9/5RRzsOgaK21HoHj4/1cmRjEpuxq7H+LSvKNh/fi6tsBmH
IhhLOSROIIzqH0OkZxlACh/h58mCU9RyAJmGUWWa065/rHUJcaE3pdzuQl6kV4LJ
XdT4G1R7ktNthku3fDtyjoKkIY65yJ4g78ukoqn4yoA0a816kal+hVnIfjpmt7Mm
Lx7SgQ8cdMiSvQ9O5K8VSJOyGoWrPPasRWi2/x87/hp7xAXNP+ke1t3aiAGbuGUe
/J0KlLb4YleRN0zah7fHy8d/Us229k0f9iS6CnruyTm1ZdZHZK+QQ0wsRMGwUe5c
nzEBdgMxEt4kSpiwhoahdTx4dkwksUeSNAx53FulWW6pqE/6ZaNCniLSy3HaXSCL
KDgCLwpQPVDrzJHRJ1nDfBBy/kw//IGjXF6kRnBhhwd4d03svbiMu9HkDWnmvpAO
OoHZWLOFkrJ6pRrAam81jFXp8hHYX4tLrY9ksItA3KXKZ8FgaXs5Dr+YEPl7YhRj
7a/APAkv16GgyMRmTFTN1IZdJrc2pDsrAypRwbNTds1Tj94rc5TfDktpnr75n42P
tkaij6ARhOleh1s6njIgwZojPd9cwnOKRJrTLfrTIkwZFLW19honGjSWiZ9glBpF
M7k0InAzpq1UNuRYyv/IIqoUbt7wWcruHdcBX9WC81YHtelloqf0WoxoYEjPtY75
tqwjyFLNEK9Toh7GVXHRYaxeVVB2G37LP6QKIiwJQejFNNBfnZv5b5MTAxcVJOTc
S2x/UvaOSubbAzJmUUFota6GQibKtrUZSXqDaJV120ryxWaMQrY+ySyNv4/Nf4X3
IfDmUzmb/P28FgQuZ0Ba4sS7TVMOWP9Ka1zRZPqBjEgY/fsfT8Rq0LbMRQGVXqrf
Pu97v6li7+YWJ5o7kM8A6n02NPX6sQxvZgVmbVdkVk46FehzQPHR3pvYroMsIROm
/RzaZY/0gJAgTk7+Ay458meS2nO7F2mTvMcpcxNybc0/RJrWvCbhpRQzYA7KsTvb
f/xuOGgMYpQO+mSBQ0YeK84IGQF6EqtxX/UDhmNKbozKWZgRaec8MJplZ1VDG//f
cV+/KfBWvFZeYRFjB/MGcWA+hp3T1CNXHu/CJkTnZAWlHk0Q9aKBHbE3qJfHKKA0
mdvtcjyZjEvNK2OsT0j/QbhGylByQwROIORkO9cK9BzM0epANssUbuXALA7aeusO
4fRNIgwhf2NRxyn25TMocyaIUiC/KTRuUUkGgR8zXmTHx8h8o8hrjhvomVTLnKpH
56erNlAKk25Shs4D6XpRYf3MwbmXTzbP3eWdxo8seHWZtHVFfZE5icBeKJM0Aqty
bgOp6QE5rVD91hBCjOnrllyhizToMtzqzenxCokRwECm5y2ahPSGLAfPFKsTMdb8
TWn6FpbdRtLTBp2CxF8QvYCVqC2lf6XyMgqWstBm5/P2ZTj+s1ivT3rnibzTN/g/
jQus/DqzJZrPYyCr5rW0SmQ47l59v3igiIfvnGh9bE4iPy7TsPgFY/ufN+90ZeEc
UI5SDMy3oYOisRpgmb2tT+d58/S2l41ngUMktaOj7hZnHmj+dpOgbIh1LKo5awns
G2JNhGqG9K2bmeEbDPHgPi9182zb9KOGhTqJi5I1PRNp/RpxbdaZclN1aK5oa4nF
UCxaDNU0zZ1gs5bd1BC4821V7V54XKQSC+zx78IhGjdPQU1VZdnNewTw6xiKluav
ncV3ZC3TRHA48MyeJ30IcMFGRaRW1ES/UBV0JAdbikHUhHGcsDLOJ/rwGqbQ2+pP
q87515+KVSIRw9hbpqBNBO9xCBlDP3yeEcG2qXmxu5RN5KHn0RxW5Ljn+X4Jw3yp
br+fPJFsb/c1fvnyDFWSLJa8Ph4Mbo3+fy/5KKgV3GttVDBJjq2S6S1H2tALCc4h
C8yNK8HydAjYE+cCCyb7NSxL6AgLbmCscHEdQbxT0Oiz4bFun0jNSOYesTQXL3oC
C5MJiOSAWKzp0VYpA/eQui3A/R+1NpccPK3xTp8WIHrMX5iTRExwkaQMqbn70dwM
4amMMD8ydbnJ0YgTpkctSb3tx3BeIsy3owI0WCdsReqT3/RZFbI7Uruh0DICFLK/
fo6sECVQn85X7Q9y4BFYwQ2J3r1Ygl1k3vHVOK2ccCSBDJoSVlNrhqNozqfHG3Vg
7/CoSm/MUaNUhHjL0tmqStFENLsMO1wr5gc+wcTRH26Dny7ASIpoDPL9on1KTfek
Pbvt6sFI6YoAtvpncjnUISrPToUqBl50V/PUkdLK6ZWo99WuSt0I7BjaYMKPLiGL
Zim+zr2U1lgi/2F9fnwZ0EWD+6l+uYH2u/DgFKVzA/RSQYW1Mce5om2xsRvL3kiP
BgcJvbctMQafLAjE35r6U/3+0EIWDgLhfHN9d8bCERvuouBXNusRS0JfrTf/j09D
Lqg9rS0x5aX3I78RzElk9m6rm60gp/KzqZWER5sYtkXzzq7UQH4pT+S4zTxR3fvh
jdaxNUnIAYl+ws0BDVehoL2akldZwQVPUy5LQr8QZfJj5NfKxHFLs4ZYGdhCxnNf
iwigPDf32MxIPoGCZzjb/X0Ov1Leww1BGh16/9aw4eM/HLYVSptKlT/v9hPMThd5
UuJlc1DvsnAeMUyBnG65EXvpVZV3CBgDSxIvu03NFEcwe02B2DjWAV/2QWe0WIpx
GL7wGKvpY8EJlQuHxlyqUDTmvRJfR0cG2nCb1T4XSFe5NU+ldQqSfSbFAg/NOOQe
thjvf6rAP5QfOFefEpg3jlHN/xQzojsny6RIR3i3+zorkOjcKVgS1SxLoCHefgrx
JzCJ/3WfIWMS87u6Us4Sau/j+hrJ5pbNKq8mHaZo0D/tzIG1J9EpkENHiAAYuIzn
sPtfxrIgCZAPxGt0xo02CDMYWrqW8dsKrEmU7xZEmZs3AEf8cDvZLryfrc/7jy68
8Y1pL9GoBJygZHZ2BO4LGHzIUlVMGfQlV2h5oqMMBuO3dzck1qR8+g4ttcIdprYi
WRbjl9z6QKOp+ffpMxFkjPFvPIibGzs2yul4Pl8Ulp+dizXeZkPHTqO3KUC+C+tC
SAPNr/8Rt+JdVSA4UlDoPNCYCM6JaSmC8wSmAVda0o/yAOPY8JapRbZ3XYTQkznB
aDDsKY4BZm1WuVQxh2vcQqMjSpuTH5l01EwkbVcCrwliILkfOWJ4SdvFSez3krS5
ovgCF0RtJfpXxQc/LrwCPWAbVvU+rKo4w+94WCYm2GsWhxTllr4hhiMy0aeROblM
gFeQuZT2YM49pUr+ZdTxLzchAyWdFu0gVj5jU9vQ6GNP7FVrgo9ud7YpLfHBOirr
5yd2cg6TGPGhWtLRTt0yMTNZHk1Gj71SdjtiCgaetp+TAKOtpwIUI9OaECRdOQ7p
RWZ9qQJs16zBytvA9a7NgoSBgp+yx26AtQXhQ6ErUgtHbXVT4TuJJ2DBGyyFJTCO
RWHMePwF5xrPjHB1ZoUuA8DOvynCALZtNzy3RD9o2c+CzRGwnUMddSCQbKrnaMoR
567ul7XmrpisnrwbQLFwh27/5JoDVn6OjRm+/C/FMykoE1nt/jAnSUMVbxAjyvKB
Qc4g+2pfdLD3wKfBH2kuWShtK17OxdStA0ynhuAEZfThl3WpfMhXTly/a6uocHMU
7EitWr4BUe2qDlK3ZwQ/0PZKX+5Jt5lmWTYL2PrHhZrxsmE82GSJBVeJRGK8UkM/
rJZCjLcczqcxifC9bXQ29FY0wqaHpjMldqqLZ2XKo6wUX/my6Mr859dQB7cWfN2D
KuAy5m7DYxzHqbMihSnzZOEX0ba5g6+GPGMbwa4CzhoY8PMCuLUPvO9CQ0yrTqNK
qpBCsNAaRC92Ob8ZrmIwBq2YqnwmWkVNL8IwxpN0r4+0HwstTTi2+PX40fZa5pjv
Ndze2oPufdgr4ajBEm8vRJymvhjrNkZw8N9mXY4KQQJKwaDPBMQdFV1eiZ/gOWdJ
M3pxCnb/zNiqfdB3Q3OjAO4ZvBwHgm+2HWtv5wGYzZF7BvFg6DhxEekQl9DQWXrK
5tEVM1RdQT+9hj8v3EGcwyWykAQ7AgODzldiJ3KSFBit8QxLYBZzdFw8cIYxKCgI
zS5BrvwDCSRZ2VdYirMvYOLIr/JH613BbWNewm8tbePBNgJDmiC9bdUyISu+QP83
WOtl79wW/h01bPoYIgmApil2H2ayx2KFvKPx1xwv6hLc46Dkd33IUmKbi7ToiJvH
6ywwNJ1jHeX1rrm/8cTSBAfigip9zBtv5dCrAJ7yuDeEujNkpnuKTzXwKDGd2RgY
yj7+1kMxmi2JtGEWgLJzwdxCoPkVNSavmUHwpfc5SfRYBAr8PgF2J4R7W2KqQCJ+
dbS/StikFYZOtBfuaVFb73Ko/EI5YtENdWKN9BaqsRs4llhjIo2yqW79vKMBLQMn
0jraWx3MmLDCXHeZGEy7z4a7+TLQ42Ghk4uxjr3qp1WnJEG+Ctga/J1ytEvcbBvw
jdO0PyKc63Dp3ToaSjbJ1s/QbQXD+r09tY6mWgPemhkbGwWXPsPiPi5HSASBa/aY
uw0ouneCncJowUrhl23lygscnOdrvNirYIryqiDxxwCOmSj2+VPjS+CBKXyq7cUB
7Nk6qKfXl/plHZaHMynNXbtGTq0vBk0RuIE0E4j8aZl8gRcJmgzF8uhWW3mfOV8a
BxgoHU8m71L9U52lUHWHRnQJgXmF/z39EmeK8ZzZ59lMVyvIeeZcvtyKg/mSZswM
mYk9ez3myxt2Gphpsd8uGPrzC9gXMYcG6jO3Jrra4HfF6jSNyqDK2S9mpNDK8P5F
HN/xLn4wT2Pd9G+dIHonZnYc8emNwdfSCnABJY/Ed94T8vd2D4+2/xmR8jYtKQPU
Xs9A6IYRQeOFyPOTz9em1egInoUs6JUAdfSY35PTyGXgwTmJJwg4FvlG0aZAq1ms
yqcnLkyBsbZ3h67/gyqpjZCJ1mn1i03+d0Zkl8ajr58+34f+OahDGhRLaj/h1QuP
Qc8qfEXXAETiYpPbC6+2AgPhckghFd0Gtegt7dye4B3sCGhdr7+sHsCbGLV+Bswb
skiY8i/2IJc7KwWDS5frS+DJfs3kJEqj6JsrSB9Ic+OFvz8SrX5ceAZ7X4X0UYdY
2hZHrNG/12XjBgv9dZtr4kyjjDgzNQJJ4WRqAUGE+jzf8L5VcVeGoRC6E6NJaQja
H2KuaYTgP/n/7r10TODpaXFTLANx7QriYqngND3hsog4JHt6CZKhxQRTNXyrYvWB
gFYCwGijR8vZ0z/qynEvjQje1OWBCIEAhsVZ7VWnD8DyYDx6oqwlaCnYo6S15E/U
YGEtx2hDlKfV3NyisJtkYwL69UFc9wkr6ANzhDQukQd6yx2sB2OAr6rKPzHh/lPh
l5+zeQ2Rgqm3Yr0y9L+O4ZpWnHhvMLoTtBumQa4dKiMAy8csFxEIVVQPeq36ZKbT
OpUbSwG2EypNtIgjq4tErpJ5enKDHNxA1i/rHsM7yHoDdp6KMj4cS/qf5PKxShMN
e7Oo3qZRchJNwLBV4DxQto9oGky69zICXxnTszSNGm5fHm1dmkx76EV//U2Ce0dT
5+misC9CIocChvxbso3hLDaXS4ObSwbSW0Dxt30tD9HzlIUf2Ga5wRQZWGucUhsy
WKFpZKeANA1HfoE4lH9U0FWFPvhyDV2NXo3nvJvNEWpMQeUG7bhUmU/BG2sTj7KT
3rfNSVzrFVCokKLD17UyfNvO6JmvzW1OuWAhjLlHXCHZeOisSBDa5m2Aehwhg24W
G/tuLfMNj8mY/txOkb1fHaavg/7+YgtlRnrf4aIr7za/MDvIwxqmgIQdIkFFnOSu
iBG6fwUQoaXLnz9m84KXLcp6+iKWWxJ+S4M3ipmCmVC/vMgmFqHCLMuMBYGFwR6p
iAwA4TSY5rtUq4C3DE2vxjGBg1E/Sr43cHXCBb2biyXh78WEAJKktxSNk1b/fhrp
OkdLTtMF+jmhCwThA2oZ90GpunJVFV1hV7oUzLL0Ux1Wv3yytv39mdyvR3fvH6nv
Pj2WEBWgRNwVmTwRv7X+iVDSLL1JBqzk/iSthVNW5bbV3xrkox2b/f5V0w51SEv8
o+WtxBgeUulgzWpM123qEIJCSaeXqEpzz8NWIPBZu+9cou7BUy8mUwfZhabab/tC
vJsfeLt6BOwWrz1isjQp6rOyLmrwhOrvftEjSaFgQFiCS+wLKEWnvYtKnhPjUER/
YogtD7NbhXW/Uc030yc5/cGWvLyTd2QCPbEZ3UIzrtAPkEDd22GVSzWt+ELGCdfx
U8WXILbWrlmIpwPe7fY4WVarexElaLVun4Cl1vpTGx27BjhJC/t6DlrHKpDPLH63
CEetfL6FtaWkK2eO+n9qX5U1j7ZMUwLAz36g0ZR0MaL2brtZrA78vgKZZAOs4GZe
bQZk45v/e7WlXxX1zpxJwG0MlMap+eNZ2VjV50JJp/CIIxmTHbCto5Vvw6Og73gq
WLc2uQQyXEIOw5UV0/G6EAgARikgwf+GVVxgDVeLBOy2+Ot9uOiwv2KyDYtbZfiG
oh5aBJXXL5LnHGGKD+6LP09evXVK86lpFtNoofarKVIE+jXGBjEvL3ezB2C2AWKZ
jK4ismRmzvCaLtU28mtXlA4KK+pqlH8peYdKuGvShqeCPP8q3NmxGEbM3g87UPHg
Z++43NX4F42k/D499L7Ets52pxs2vtCvelvPDolQ+laGaqDP0gJ4PbBRKDHoyu5m
ImrqWBQa9asBFV62mSOyyTniaFl8CV5Tuk8WsAC2EfA6RT8zFWxtgkm9BPswzYK3
E8SlTedvi44hPd3dqv+21O3WkMwRKu7XqB0VdZUu+AFqQ8wseilKtN9rzU8JCA9z
TYttV4A6vKZYASm9Nm6OrAYdYC+9h5uM+H/kmR8jwrPpS6rov0b9oPbg5E8idkKh
LDRKlLRTbP89eQWcGhtRscYTaI49E2R21czOUWgttT8cRaZucnSxksJtow5Vsnym
2zgJTvUsz+CHWhHlsfH4aGjTK3Sj4CQMv/r3iGRAp9Sa7o+3jhbRn5fETDdm65Ch
LwRx8HlgcRjvBwGvmbo/OnQlrSV/2p0ERIynbrNVssWErqXzuHBNixgDc4lLe0By
sbFBz/TsGEzsTcRwwNd9DKK8ogIgCbKgxgXwQkzLgWNTpb6/K+3WoAgVuVkCnsBN
WvYvbpi6+oWoHbxs9LEbv4Fa+OHJAivnWbcoGYpByN57bYsFPmvIYI1e5HqJDtCV
3TGmWyRGVZdzrDLAUJ7DXn2Mdcz7PUs1DZXEyf3NPHgTeZpKmFRto8ttbIc9hrk8
seaHIO79vBiG5dkpmr7bcpc5sRtUyM0McP1nBj/vTIfkU1PS4aAOd4/M38o8Rh5Q
wi//hX/120jyVf5hfRott+S6gDhOKYfsjmF6Bs7UpbMLeumy3kgeWBZMB10DFvgk
8+4QVUWg9sHOu3aNYu4J0k/Vr2eryIVZVhmViPfq7CqHbqa7qz64J09m3aKLfilG
+doVbbzv0WRg44HMfjZgLdYihL61i+bL86zQKNtD6HxXycanADMqXAa4fHbZVdJv
Ox6B/q8y71Hc9qUj9h6rC/Oiqe45CGe7rH3qHXINJPvPofCqyh/yKgORku0IDvoU
4onNG6HmGGyX5NpfIikbR/TFZe3wUYG8B7vObNOuKLPsM7Zn7nG4dhieKLungMt+
Wwo126NSbpDT2BMm8LCEim236YPbwODcVHfSD9W24VktttyQ9X6GuqGcn0KblCgj
xqLOdL0yXKAP+u9j23AURcsAHkJrJCqf5SbyjIlmSQZyy+app7V5+JS52WuHGh0r
zfp3CghodTUysJVJeiAEKnd87iCztA0EvJU1lyz2uBswt0eaxFsPYW/nYRUh4YX6
S9elPubJ2FIRorni8bjW+cmGa4xqDvL8yTyNsQAK9INm8z0s3CFXIwlmpbN348bh
h3TfKZdN3kIOzbcgBlzrFWlvkcoKiEjQYq0RgB/7D8gm/CThJVRoJWOCJkRl+zJ+
8q4GojEep+lyg4ba3CmntdBxqZO+gGBWVLb0BNuY44/eGJIsZ7Ki1+GVS2gGK/ML
1li2+py4+1ecLWRQ76Ojm/AU40eMlqAyAeDOveflWI6s6KwsJdVnB54AfH3I7RZC
Bp8DA2uKW7stv1CHjS8vwAXR4xQuZJL5oX32H6o8d6lL2inhb6Lok+CUf9Wr1Koz
AL5g2Rwz1GbimCB5fjMVcauwOoP8BSuAeRRW5g3Zd+ic+Y61XAnrDmDLFVq3Gm/w
L24Q/O/9Y3Bx7PA2t0Is/6xG8+5adXE2+hHl+5BV2tX0q2Nl60p1BpZCh5xSuwDS
r8ctiVm0Hm8VNmEso5dkEEKtPhtESqwx2M1qj9dAJGHkXfeQanTCx/sbgTjx4gxU
LBYoxGgwFyvLhxoWvOtwJ4SrLX/PTYO8eLd7YXB/t5Q/ZGEvkzdCJVoU1N+CNqVh
gp3MTP1AbZwDDESgVQYssMmkhOZcOrJL7tlb6awNEahThjHxDziBa9gbYAm/QzY2
4OJH9nvOG4xwDCaODYgvgtfzu4VRr0XApvf7/Jt3Z0iCRgM0TOzLp3BvYfChEUok
5SwRowYUrIQw29pHggpQ2LV0j8n4bk0yRqPDH7h5bABC9qv/ScNUdcrgQK0cXEKJ
nXHsw99zyrA9ZOxzMs3AsJYZHclc3e3vyTJwsmTCU5VDs+VtaW4FL+Mh3cIBYX3T
vtPvRA2LrcRqrYZoANQfO1X1ifx2NPjf/cE6rFGumdcgONLJZhMpjEurZ0bVZGOk
K2suH/EYp1pGYO+FCeiuSln60f9CQ3QeLe8LLqerjeV5PQ3Oyr/xodYMU26QLg0g
6/07SWLrnMAMXC50yu7yOr+u6iFN3t8tazbi+Ya6qtDBh+mzvQL47LcBxHVKGO1t
1c2rBgLiTwc2E7vRO9spqOh5Wddk19mt/s0gMNCl9Uxdncovvu4SpCBKo+9TSQNh
qya5M4Wzh1DLXz8odlxrdVq+ZqaVFevOdzh+CTXzzwLl/tzyVDPK2q9Gvmze3Aol
MjhGMPIA/QIe4B+l5tBu+X7xBISgCrE+k9qYjlCihKNG6k9Yw39PYZjr7VNHfbzE
rg+FhrYSUJmcfpvMQ59qDJb6zsR2ONmF5R/IAPYefKM2nrLPuseRbtNkDqxA1yVy
6d2xFSHh236gP3l6pwkGE5ctzFZdEH0ZDq9/oLX0W4yG9lBmXKb6AV429cKDYk5i
BaQNmSPcV1m4dZ1zb4QYbGmySapkWYlkMxsykbgAc91uYbFrREZu1aIybwI5RyKK
PLSjzajRbx94OFRbdkD9Ao7wIhFd/d/fgQzwpGQ4LHAo150oytikXVk8YROn7djo
eJ8JMJeexuGbv033VjzTud3LDe1PqikEnyXgCCGDmVAFU5i7dpr/14Cc5lKDpd/W
GjH0Vcdrwts7SiRS20NphEePS3mAeUFdVE2q/Erd+74eoEeElJgnuABfRgj/lNag
rBBNiYFmJABa9ervrgVALnBjg+WHIThxoce+NtkxrCUIddxB/RnEyVm1z31xyjc8
8NjIGIyngp5qqxj+6mDu6ierevsu9FkVhjJ7AbePBWxKSQkDa2DS/KN2FzuvEJat
cWK01xD0jWAgpaccC4tkFIIxBqaHN4W/OOFB7fMZH938JsB4bvFYB2oLVmHEiSVK
T8GvWj+jbvGkizeeFWiuAUlsp0nC29QRMHx/XBTxzUTHtFE1wURJ0G34ivGcvTW3
xCszHb2JE3+eLryUQMja51rI7PinTrIhLM5FMOOjZ9FnvkhsqAlPYbEeClFa2+s9
9vE3LqMy5MCWWCkZptl+amPkuxIWvmsvAhNklO3Vysd3NZGJtlZyWYWy08CmjKMS
K92ork6lx1IXjsEfhSkHPuCWQEY7c5prEYcpbW2h/joKKhM1c7Rszw/6zAd2uTcI
5dDHQJpPcD5gZf6rI8nXdwjB2iWHuEEMvHI+ODe+DG3j6Ej7xNuOc2HYFRSZu8FM
kkq0Aa59Xg8Js/0qfwOCFF8uyLCsFkFeu0sIG2+LWeEdbnLcMifSoqsX2RF+XeAs
xUfticulUyjBzrcyH6DwaYRl3FKLBcCIu0rOgOQFUv6GBAaJtFaT7aw1v//sxeRK
uRQCxbrpw6LqheAc9kpfhDf21RuwA8sol86gQNsITLCd5B0hz5sXZLYsQfN2Cgct
GEA7L1Z/+xpLUd/MdVuJ7skounOHO/3MDCY8L6bc1cDKNOyp0TOuPfO8Jy2bECM1
mW/KYCrWElQWwD+aCjGBYSPO6GTmjpyblGS05k6mR1NFWRiYOOvizLAb2taSxFOw
YDnSFznWMbdITTB6hCb46I2n2bn7Oo3w+YmGpmVx7VGkwdpg6BCVa3ClJZCFhM5g
j3oxkGHqYOUnUZcKNpH1lV5nHxLCuFuwbbHSsFen6wT/mCwdWNZ2YQkdkEedF1QL
Y9gI3EHD4O7pzX9kzeGEWjT5myLDS/2n5wA07ztQcApbFaceD9XXaapG5Y0ak/GA
6ssS+mMAOMlW6O/W0OPl96ATmzsjXQvx9BuJuH68sQYRKSbtvKkYSDTXRkp4hERK
RVWHw745vg6QwgDyQ2Sg6Pn709Wuo3wC0IkCVDdgDMXUCa2bLLiF56/F/fpqvK/V
5PFTK+ItosTGD9PzAKmdNyNIRCv/4qT1W/Y2SkA5hkR4kHEr82cut2I7u7QJbO4k
lsRdcUhgEjumJ+8QR4S+OuBWCfp2h3wYZq3IyC4MHxLqPDZbYxGZTIZFhSZkPurm
vofv16T1xsMkwVt/c5Vp5XbvwU4mPRYoqxB411v5U1UA9Nvqwm0BmXwaxOZLaLPG
e9795kQ9JDwl7Uvs0OVvlm7B1pm3UIXAoDBUzTOK3CPp3WAMbcXAzv7PpxPCSjX+
afIjUTH2i1yZTsFpml6Z82Ol38rCG1lgs3Wk+aICPQO3jd3gd9dn/B/7zEVhYYMC
F7/emazQDNe20ke0t274xGWkthlY++oHbs7bbQojBnOvYc9HfdqUf1zeUhN/EwWm
BdeQYITJM8QiOVfilKco/nP1KeAN+JmwSEqk7VpTPO0U/1csmJus0NHHBhnZ4JW4
xbs8neYBqI/fOUzc6gTi0xJhSxDp5hMFhWCgDzfwsaWqBFw4vWNX9gAhgEqm+v+Z
gjmb07G2JDqHZV/ellUoSKvQZmFeZWaI2JsCFNj4RpEMpdoFrD5VqvjfUTdG1hrl
uaiDQ8P4ID9wC58jEIT3E7VWcmzxKfgaldTFJ0kTbztiNXId9+s7806FuG6jtIev
4VJPbZgl+qdh1Q9zzii+RL35ypFfVAM3nAe2Kq+O4dH69yWbTNyik+OP2Rf+JCo6
1DMIISHew/evoHNrzIYIUhgbJaRzpcSmqh73/DXs8tLDwt85B8f8QSz+qJzffrWN
wDZ371RUIGq7ziomh9SBCVBi8JuCqQrKaYh2I5wsCWKK+ZMBqnxgimqNjspX9JQc
fnal64bbONu8R/JRmeeJPJCSQ5jWZVJxZDunuoT8hz7Jl48SGvQft5LyfuxKtAU3
pgf0hRxUu3bKHqqnz1nTEuWzR9H40ipX3DkQpiMxAWAf8gNVrLpjXJSfBJb2MruF
q9tT2PMnu6B7SgZebpExcFT2szekiItXR/CaiwjxDdzOlh7UjQ/Ompvdr/6lu/mX
WefiIzUU668yuF0cE8wJ1Kbp6OjOfgdy1IXF317N3bLGCwqTMaQfnM6J5Eaymgnh
n73xdSqbd21zFsdes/d/ahQJ4G0EMUD45DBQcd6RN0AQs68g4EzSo+LVPF0lnAF8
XMGZBzHMgSLhPNsgtCTz8StdjuZ7jSvi47HA2IcRR9ZN37mIzmoGAcEJ/aM5kdjR
VyTbBJ9a3NSr25ykeb/VdYBD6bAtvV9QgX6df5+H7ntbxJX/sNvl/XjfXu8LZa2L
F7HwD7US2uKECbtis5rhwe3ch0cwwki6017lcJFR0sxqqbetn4rORQ2YO+OojXnw
UC7zKrHMgCTdxfVSAuxGNYAjkbCRYUggZIICP3ZNKAbqPKxa77uIVLy4qK2Va6gB
EpGLKiGgJEEoUAyQiZ/oSCWiZ+aytR1anzahj3pg63kzoULGWY1wKA13ea70yNH4
NYeWwcZjNmQaq9iSzcgaxpAx5SyVbs0ZSbqY8mRZcuCxdHSJrFaaL237EUwUiOLB
mqo9R9mV41eN46etvHl/Y0JBg0a1VEd5N5BbIFEjFYGeEEySrqzuwhZ8ZPd8GZXi
3O7kqbEOojCdZdnAc82lgwL3CUBrU9d/0k3oDY6h9113bw1cIkmb0XSH2G2uWeue
HfRjGAWMjJmbPdoEzWfaE0jrcWcbkqcoUJoOoRTAMYhaM4g0EhS0UoGe7H6FEYYR
rb/X4JCDO+8Dtu95d3ayP52H8v63m5X0vuaS+pnwOjWv2zCohAt4bwG288/xKiwm
82asObHNCuQxjDrXfPk3RaMNDn4F1FV43zl+8oUhuuuyJ/xdpvT45L8YfcKcxrG0
4qs6tqM0bjqKWJTOqA8abpG7ZevmKmwTZzxTF67Ap5Lkbu3RYmW2iWjScKu7+FOQ
fwm4g1GwuzTzrdqSC6L7lo11napUVmeOxtS/oeKOWI+Zn/P/mExZSpbAtkItwrsJ
FvD4Ee7glysDh6mMhpZl5A0/ir3JWaUeWRKhfbSrS0gIpYFnCO7iQXUXZowySUZe
5D3XVZx9lSEcN07ZH4iH7SQyklPQTfFjaYNMm5MN2JgBDXYlo7/oPFWvgMOk59BQ
AoLkZpk8Pcz+ph1URCLC6z9sCbQC1rFT25IyX6P/CUEqA1pHhJEhMJ7ZcrjpjsJa
BMLUFeRkpFnO5uMXdtgHRBOZ2XaYdHPXgOcZHeROU6IkbdprqOl3jJ5bVOLWREtJ
TTTMTsBqa0UuWFVYL5XkoySBjKhh3NNNnzM2jZHJG4o8QW16AWs79Ibjma0TabrM
UIhplA4VUOgt/NMTGPIte2imwGZT8ibB02dMpzLihKF2RITrHyrTBuqlNcwo9hNI
B1JcFHqh6dYqOrfWotrg2MaE8BAS2Icqd0BkttLoqmQwesin9TYcEWyaQV+eM4y9
KigIPQdDSwJZuo3Zb9O6xYHYL/FKhFf9QpLZ401LjsASnBIsk9ThCwmvoEullV1B
WrHdU35GJYSvhKfNeYO7h4OPYmo9VCu5/F4kLkRu3Po8KLYZ90LgKE1Jn296i5Nx
mZc6ZfYvtCq8aK15vKk+alXFYfUWpTDkBbYwB1SLhXPTmPOEo4bGet3HEWor88CB
uWbrvn00CcK+mLin8N9nAI74SC4fT89WLtJbcJL2jc/bZVqNm/JYXQAHG7ztSxE7
57/6LV2PmIZcMWYcshFUwf7BGse35GLwsB/Iynf5PpettK1T5dgmjN5QUriBGrUT
g/6c+jHd/4v4ahYBjMvnDSTO7HKzCPPqFtYGzh8qtY6JOrDUZMlH4pK5Gaxc3zZ+
R+XOW2M+MfVhxaBtSyDTCnZxZ2OKthZV1F/FLyfPxAcolAdtnHxlRMQtezGB6Qrz
d9gxdJkUMsBXAg+jvTSjlobvrVgFjQGBcF8KbPPNG5MGRQddr7i39Ara057FUtaE
WBK8AW3B8j0KQJqai69vpZolUS4Zl24sD7x8BWUUR8zocDunRJUk/7t+GhC/8DfM
Qu1LGRYgUvoa/wtHuAHOpXUiLuhoSKNtkFl6sw9FVJsHPOz15Cr72wa/O6ODYr0X
ZDTJz1e20zKFOvLbhgqEVHBVM2QT9zR1bvKZwqbcNf5zPo1TXjFj6fO1uJy0oFg+
KbwiMHWKKqnERfMyNV/XkZvm6J4Hf66iDw2fc4OhzqkhZ5TicR9QRtOC6ozs3/We
uoQVDJCmrQ5kC50qjTKer95wmQtaUmaRin+Hk9+QP6iovhFdV/IMV4lVniocWunQ
Fpa9PEiwRUbUiI9+R/VIBUqzhdEENiUgbFI/tpYCoaUYOHBdctQ67I4bbi/3l/9a
VIk5EtDA+qfLGVzT0Jnt7BPhWeOcBYuYekWF9wHmNwdRPYwD2Ii45C5nUJw3kNrm
MDsc8RGK10r4fPJG24b+hYp2IvTUdl7CE8v1z5rNrZmJDhooU9KUkYhXWg3XP/nL
6nJhvKKT8SpO/oa2UKnA5nHFEUbF7tJb6y1wlUC+/hJh4jw91PMXBtWbQcQpcgR3
q/XU8BpeSbHa6gFsiyWG/pjFOXwmiOljTGmavy6WfphnKEy7V6pyYY/IgPDrZGwY
vjqSn7P6b7f3MS+tyvqmZs/9t4Ez1x7ehGAvJuF9Jqp5lNxMmaoOI9Hmu2/FVxm5
9nijo4mPzDsEr298pq1+Y3xC3l+bjQ9H5vXbrF90GJxnL5UsTX0NcXanz7ZkDJ6s
yKnYMeW6VtsAT9bYFN7un/ynZeF5ElenwYinwAv7RyvBnFu4X9S5y8rPF+kWCXjY
XC3rsTHz3DgTU5B3ol1vDG9NEMfCJeL4QdQLIidsEmPzJ9TJVYAUqarN7bicY4fc
1LER5PpUcD7DhtafWGv6T8081QdIi7zfLSInbJB23Juyo9NZ51j/C3N/YBarKpe2
LtimdhXw6Z85/Mnf627jtraihsxJo3+ik8UIfGAY1Q1THDM0IDJnFyc1Jt6g096x
Ne89meUmE4GPRXS73VcvFluKzonU2gJHO3++WE/916d2cEIcrkS0pE6BH04SXNRO
ToUzG+M3R0mzs2m2YIsJJADDyE+Pf6G2cc4xkh4uRVoeBYnsuWl9bn9Wgrn8Nn9u
t+VXFcVj7l7TK9CX9ojQLuGBMTWRL7IDA9MxDMxYGlG5JnSWt7f+Vdm3Lec/9owd
lo9BkBKJEHHycw1JtX/9UC24uLtWffophufBX2zsuMy+JL8buh77o4cyPCxRzLf+
bM8HIt2BBvN8RV5z1hS251SVLu4nkkYFp7uRYCIpsvLkNrXm5yYuqg6dcm+pdmEP
PaR1f0/OFB/hSzzKopJ/wZwcIy5xd9xz446vwExdT9jAAXhZL6VWiJa2A39/M+MK
zu/vFlQxzZki4lXnvX0OY3nV8AL8oF9CdKvOAAV8brvVwnzbgjFjnl13/OJp52tC
QlqfxC9E5wMeLHPGa9DmXfWTWoSyfqiJBaPRC7ksh2Y/8Q/B4G2Gg7nh2PrW+hOM
1FSlnykx0RY1Vq2Boq+fOaNrMrpPB5W6POl8KhhrbQ9KYkdMw6ni3iweVZgH8/PQ
5ONnHnvHpJLPVRyMSHTGPsIyRFaGOi4zXV6oatUig55J2pJm+Nef/QNhe3z4R+yd
pe7x7+3i9ZAntL8Wyzz+6OTnP6lSDl+XkTV+O1vC2bU+Iov57xAJL9uI24n+ZumA
/vM17ujjA4L+ZyR1C6rZHzzGzXdvIthkKtYGiQcqxRkCS9P/3B/En2qm+R2K3iZJ
Zvt2/ptF+O01lpSH6x8fj8xG1fzz4s9U9gU0pvv7O24xCyU4KsNhXZl3D8gOmTHh
8LGxNX3vUcBfJSxizYWPy9fmC4GxemPnxQ7005P1GIzPk2UHE8usoPN8DUFhVW/v
WKttXOAJY7c3bzUS3MpjvIQNF2212apGar4sswKz1aEBmA1tu8gMin3S5OXFMVck
hiubIDdDzujq8GQFr9HH8nbVnInvLIAjMx5+tvHLKXeBLK0eYTR9sYeaMfC+H7sO
ipya7a08GQDhNNBYKbPo4vDr+GOhBWR9EgRFKElENmUPpo382IQRYalQEn1SvENe
9hsLU9oJv4lKMfWHWwf/rxXyiZMKHFg/pZ3tJLBiDs11S8Ny2XFF6ktyQX3nWWBT
nOMoUWxOt3Vil7R98WbZsBR5eygfpYW+E2TERT8t2CbM3pPjAajroX1n4Tt1P3ST
F+oS8TPcGzGh7XZl4dO6XPX1YoMfFhrfJ0olW2dSqqg4TjOBbHHbnskkdEs5Mk09
NOKfL47TeUFwrLmQ8DYhgD/EQ+fi/dEMBHjf9jOnjWnFdYFcrwMgH84qefDRUwnq
/5HrOfY4pfl4z+kp8LHhHDnIo6C6rdx1Ed1sAzbyFhYhBIVyX31wgAzz3bn5i8MY
ynYp6AO3t0TVqDo3KvepGTbKh8p+rJF/4MWhR4JWlMx2C1Yw1rRl4YKn5FnNuJGt
3iUEKwg//GGs6WBCz/gJy4Nb3n6t4gGT/bdBdl/I4cOuP9t/BW9+65n57OWUdiJE
0wmjRsxD5TGHt/g3s+HzJ8A1qrlJ4BjR/9iV9fG6m1lksVmVgIOpe+S91PML4WND
zCfNF1lWP8s9kL4wz8pZVSb1tw395qsp0Iu3chkHP10vkqM+NcsLxMSwoPJ6rsFx
9Ee0DepazGgPYoJsvFlX3MubWUlYYHIIhh2sZ4c6bmvj2qK7KiP2Mcdpfmv7D3Ri
vbI1Pcp+UTL7Gpo3fE4bVToJRI2huWQpzKGZb4qjSgVuZb7juwoTriFY6JCaYP41
xTCj3oOmPxMxFDUlbpt72Eu1m5PepkYKlYCtEQakrRYBb6UExuLldVSPLN0iSg0r
hcONmfOTLe90AHNgM2Jxti+Cfhd6j5CLRlLJDV3QDBHgHdhOJ3YTXCNgc0JODzLp
ZcRQAjFK1/sCo6dHqptYpPyzjIPyjq2W66ppAWMGWe49f/z6zbwyByGp/WGtIPuS
I4QKn/BAASUjKiKM6wNET4dnUKEFmbLCrg/TTbaZ9hi1QhoMbC+sfkJlBWL9BbBM
Z+4p5fhxBXF+nJgDl4i95PzVThBcURdYOwTQVlOxPdsmY+UHk5qgcvzEjYSiYB76
wtKkQUD+Rjpk/Ql/AjFjuH2OUMF474eRRUs4Cw+8RZ+EY2RXNqiEHZcSt3O/0Kke
IqMFkBFdQy5pDmkFMwaNSL7Rs/XK7pR/Kkf6uaFftgbiEEjNGgOEGJ2eBK1LQm5N
J1dUmadJQoYhMINyTQNOE4sESVdmarY1SA+A2ce7Z+HktgoOGn6/PKZ3RjkZqjyU
7mEthpE4qQRJoNGJKBEW6Dl3HBlV//qdvA2IAfMPC71iRwJaHR0Tu4qHKrhlrlwE
PqCn9P79cO9rs/Omft7lHcndY95Aj/+/rOD/YOuS2JV69KjQXCsg21Z1onrcQja2
yx0aPkQNTg0FQL+zihz6fi+bnxtPDglVuO1DC2j6P6UYP5KOM1eGfhlTspwuL3CP
8+ehYKY6hH/t9JtZHpucjPVMAfTlBc+HWOLmzh1j/fcQuIJumx40TsxvbHXpexZ+
E2gDQrOpLSXQcznv+FjS5A4PVFQVlrNldp0dO0Z0ywRYMrXD8ehlNBO5DKYj90sZ
VJJqXs02gQwCvC2V9b7sHcmjWT+l2QQ7d9lM30/t0wosG0MjpJ7lOTlL5KhQezls
m4hUNbssQv2tTVfpCuv6vvD5BkUwUKJB+FSAy7UdUER0kNRdJZeXpnYBg6wa585B
JbohrPlT1YlMVKu3pK8os8JUQyByz6roSMDBQub3XE/VkO/J5I8sFyy0VMj6Sc3k
lZYptQizswtFS1qXj6lbIvGjt+7at3Eg5JRoTuT31sWArKPJeMM0Umn0bElwIpMs
T26M3zYYYAeu/mcyUpgJ6IQ7Qvodv/LWTuzGpNvv3KnoipdKsLvfslVexoecQi2O
S1X0fk6pQ6sHZN5NHh4Zdf2OArt7NdE0GNnFVmbksr3X60vT2jqT7+dZ8THHLJYk
5ThtPOY9unmVxer82ZuwJFISGw1RkOVPH27bmuZ19jGnU379hm43p2GNf7qAxxSv
jJVs9h5leA8jWXEifqj/Ce2tsk2c/m6aIXwMat4T28NOxICC4BM4JAO8ZbZhwmQ0
6Nm+pKc4Jh2J7I17ZkNbaqqof8TBIgeHGkn1jfB8r5Jsan5gwPXjAz/ZTwRJsKLW
BewD1kwT4HFywYRpzjimarroHXtopx4ZdSuFm3Jt+DwBPEh8tWDgI1bBaKDZMkc7
eIXJqnNFQF+LHTn6usDfUzqMKvL0YrRiM7lxc+Z7dEnac95oUNUCIhklIUlhdD2/
1EBkdrTsyRzHVrHkCKCO/fJ26X4TZyBWTdc079zwHq+zhyUjtPXwkhsYWDoAoO0u
bRQ2dta7Y3Oru7/Gftr/PLL1bOsHBvii7IDJWUrhy1ErF5B/vX4EpKobwcQn4zmM
yhIKOanl8UYqx9T3731G2usio7Q7rXpN+On8ShOjN371J6xA6fvYKBFaD/4kHeBd
Du6/HbaexK6EPaNll0RGOBxgtYIgQZc3WEa4APmUF6t5QlhNiZaF15h8aa/V2AAg
SKKfB1MjiqODxWSU4YgPWpV1Tb11/t3v9WycmHZqeI4LHLkiZ4TQQaGB5hxK76d9
cabY3wFWaJ9WQNlZe8Mm5j7VHgVdCDaxB3mKIsF2oyWvkFOV9YdNOigDkWVSfMJE
7jZarVk/53gZjyP99ntOUIZnpvSHg+56Ui6nFc79SzyyWG/MkKNUv5Ar2PLWpQjz
RiSe8mfgbzk55Gk+sTA+jFtPsKgslsbHWwOfvWaqt38SMYfB1ePiEjF9UHnMdEo0
zx3/ZKo27QVJ7zNwFmSZD5ZHuASDa/fTE15HzeYMG1XLrjjga6UEhrjj+YoRQYHn
nW4Vuqw24hKeeoK4a/Ao4bfWPcPZEQG9G0n8qADLcD9fbvOgMCw+aCPTpN9uNkvC
EbJXHppt511vku0CFZ7taETdZsElt18L0GfzW/BWKiazUQ/bmB7KmxoAnFn4YXvG
JQkdl8ZC5Qrl7w2FJeFeKkdCdmgeorreHfmGgSk6q0tQiwmpj88dK+VRf834uMCY
ylv5LLYrJm55lKRdZmtTnereF8yKAVXaYHSG1phFHz45CuanxkiS52INBcQFcAmQ
MJKKx6JY+ULPIMRvGL8r2sgFqPryRIdIbermrsTcqjy3jwYpSK25t36wKS1yP6Zd
9HZr4CGyFfmvrWucfmv5VOtaveTs1iJPsHdS9LSV+sFrlolz5nuHO8Oqw4Eu9p9r
KvZ42TX2RLkHPM1K1/UxwVXhu1xhJMc7UfEs7uWKtRD6n9xWX+jfsS9demZ+KbjQ
+xevG69ndnOufl/BMMhvKyYCS1/akpOC9/Gf4gcXCrohA2XsNf2G/yCriUIoFTgs
GzqdmXxVUDzlrsmbNFGLA50cqiMdq+QUAbcwuVEzpZi2WM6FnKZpo+P1v/OPT2Yu
UHKUZfG4JvEfsEdQWcEHJH8hLqPpDpjCHKla0crk3HqDvpjh9uoWXcL2qMn+ip0U
bSm7j7+DGHUEuJOjLnoG615/1MSTdsrgaKCZZ923pJwzmgyAvnPlXRVJABHaA2Yy
wC4vcoBYihluBOZKwPQ+NxNaQH5jTFereiI0co0ZyRG99xz/medbQ0U6nw4pNCRM
lMXZivslEhrtOGvDkJ4w7OHMF9uw7FuC/+m1e5kHWi4oRmKhSMFNS44Z2/qzdpsF
5Rn6BxtspGmOvSF0aKmYmXYwUeWMxGpoqCK8nb6iem46WPnIWrTCDIOij/LcWyX+
wPSszech1uPiEuwbvL+fbFEYbtTvhAPV7t3iOzK/0hXx9eMg1tvxDByvdVxnKmk2
9Bn7IqqFVWxW+YFb6/8ZDI+q+kHP1skypgtLZQ7LvI4aR9BX/geiCUrpzS4mSHm3
EQbkPpkHepyiwbKvXV7PX4qLOYUNdVJVOTVogL/hWXG741tyMHKmZMobkxEGLcCk
/i6JswoW3dumnIQY6hUhgfHf037MNyTUCLtLrSveV64ERLiCRw29RLCxNX5NLdij
4FZSdbH9uyfC82hdfW53WSXCc9hQJxHMUuV36chK6Hq1D9XKvDjBSN9fH0sfsMMk
Ikbfos88V9h5/PTaOeJRKRCGcFFhMxXrKAnU3QEAnyeaFK74xboGG1olPsM21wpP
6uV+MiKz1Yh8ut931gxpjUDpYRyqUcxP/RXZOhPSjrCdUDKLdUxwi60PdJ+8h1V9
yIo2hbc24i6g4G7pXutcyf/tWrutN+p4/cXaz4+4riswTa6SRgqDU0Ea1UKFdjQS
+odlEI1bA5pL7gtIru1eT/jNWACItHEBmTJcSufuAVu3wyYdpQtirrpE+S6aFBKy
y6DyuZzkVC5puBiB+AExgHGTQ1LUandinBrvSvi/804L3VheJOVlHQvwWoIzxEzv
cwlT+H/+EwV6JRu4Q3KqAgRwTg4qKEPKsHXKTp0+6R8Pfx1Ht/tNiZkNdsFZrnn9
1R8eGqP/XpdnLeNS6o2QolZJQ0BU9NkyIFrplAZXeIDXZNRAvcZUT+RAC23zoM0I
3autL+oyzkqzjzi2kQBDvWXz4pwjI724fuLHXcKJLH+6n4V8t0vtNBhQ/CvVSBYp
b1xRZJ/ZtF2cxrTe8ID/vItWS9xUGuNxpZOTKXcpNdY7ksnwCo8uiPhlfAeRAWH1
IFFjBzPwjT+O8z/VHH9zZ5JtS0nQHJcJ+/idoXu9sadY71wKHggF5xFevBOOclIX
szwm4tAp0AcOyH2WOCDPtXkhEdmrnxfLOJsbrbPaI5YjIp+5oHpjwmV+zNH2/5iP
RD4pM2SUN2LNz2NBRODVT/XEMAPhBAmyA/ubQ35uFyM09zILP9exaGNh1AJ20iSd
HkQiX8VbLmESWXGVW3WiHtb+9gZjHxE6CTR4pC0Dc4xN54pi250ZUCUo+SsyEmxE
WCfqyra4bu8fZ+f2M6HmEd7TC8lW+jpR0VRys2qSpIKsbL5UetTHHLqAVN4wtScV
vTk0vqd4z9Pmxv9vhr7io/7bLG/9Vbnn17YOXI6EaTh1GPEPAbalm/WGOgS08wOA
PGkzW/lzytwx3ZcfM5qv7J5M0Yhd1bemtBSeVtiMr8upYTlyQlJwKK//8TFK/BKG
z9c8rAZUZ2qNp93A/BuMVNAmbABydTIQHGpyCPU11/+dRjuiaAZQYdfLj37cS0S2
qN/VYnS89TAg+2iyMvSGqVQNZ+QXskgSy5xlH3g4Zbd7nERWYSukBkzzeaEhjNsG
FHaKasTUuSWctfKsME4rOf54bBe5BctLC5ALUa/2sPH0IIGAiAM6elLIvHf0858P
zNcwUnsprUSC7HLKKny8n6ZXdq5TIKQ2MKpCUxKd4D3chCR0rIDcW/Wi7lPBeNB7
GWvpOU7ymX3tGNJrB1g6P1lNAT60gmKD8S8eezmK1Gna6XJFjyi6VSpgfKoiD/4l
wSKXbt4hRGplfgG35V4OcGFu9d/KIG6Y+03HbAncV79GKQNuuCpROW0jKvKl6pvH
ranlMI9d3Jz6BZjL08RmcHCh1OLZSE0GRMZfqpfVq3gjVCCd2/zHxTttAlgT6lwl
atiLZHew4vwxqa4QHoc2/xkdiSNh0Q0bIPQYF3o+x7iPpni8a1qOQA0GuK92Btff
CFKONct8bt5p+/3iPUDjPKnVAonWIg376WZ4w6HllmzCD7rdLm8RlBYFGOweWk+q
J4Odkx5fReCsb8bcQlxl+Saq2bGkyUT3EHoQtTPeIkWV6KFpvUO5Ww9aPyqOUqzU
yiptGomI2sfiEL20PTQVapS6RAsJvmHjSqmcNzfVP6gFm1l7M4c3fJorGV81WggP
FZN8ejqJIhvUgVpuODe0ysLMLrMbqnEXD/L3MmiK2e/W/QHZDVzQDXtGn2kwUfNC
l6RAgXdDkUlRj7TZEOgabQukzmlFB790NnRVBQb+fNNGOMmjvSY0KhoDYTJsmgSO
3VU1Cz1kHjzGVWljgo8cIxw/5PyA3U58leKcvZI9h/iRzONaPB5mbFdb+w3y4ohG
0dji01tF1AwFJJ8+C0Ac/cMBIxFFiZAeEqdMlqsI9jIiGV6myVAzhJ/f4JPbFxpB
oU9xKCqAHzjD+KfMvymadSQg19V+ATwdrr9qfwlNTqW49leO9/sJ7cWlAhWXIhQl
TY5r9/6NujacnXCCz8EA2VyQhNOH3mXRnF2P+mEyGlmXaGpHmh5PbG6rsKVsT0XN
YUiljK7TC0eoCePPrWBCfY22fKu3GYjmnqEWJYC0ikpiQCylC9QxWbQ/qnfbNPmX
FztWqjrU6B3hRIKf+nm+EPuH0z63ZXsWCymjF1pWSRMvAv9h/KYM3AvuGI6SHzvR
JeTmZUZkCyY7K9O9wCKt191VLOAh0BPX6ccbKSUAgzeACt8p/ijjA5ljVIhK7mAG
wd1rlvlggrqD6uiBWKgYtAhWokCgDS+yppreEOSOydNWDVFo7/aXpSmR9ckv67mh
v3f3jlMkzK4osjhw0HV4am+atcRTVF+/ipQY5zZjHZ7fWT2cwivX+1ViowoHL6vL
dLU0YzAP1muhqAGK4GPagkWvpQKuQE/gWb3WTa9I33Z4cZy/x5xtkE8dV9MqMg7J
ZOtQO+ETvB//ctj89rDKw4+5N474CXCPdkDCsVDLBrP1QtMUGPxBussQTPvkQ5F3
QfPKkzcBLFUiNC3WaEHsAupiTn/KrbyO59uHOseJzi5maQ4IrjjPEIWH9BocN0kt
OMEZRrOm0I6pPM33lgqTwjVGKnWMakf0IOXnZ6rQt4rXBIv0F9geEqwTKWcJf00m
u5rAOdq9HgSuyk7q8jl5QVF5ytSHJ8VpEN7h+E8FYP5EaT5gp7NTJIGqRyZW1Hqp
NRhVRpZyzaNY4HZUJIDUGMG23wH3mYIxpdkDC1NgvM5XZQxb4+QfM1Y0Zp1vcz8b
DWae6eC3xQIqwl2LeNWR5ov5RtSmSaKvzS1tS5QEhR4LU46pa0LFrCPT4OMIQm4o
CTPFpZa3jFVeZAOeYaeUu880J4V8+X6h14eK3+81blVzrK/GKh+JlC6Tzd0JtZHU
PZMZ3k/PxXOA4egigxqBC+oqXxJNT8W12Jpu62TEUiqwiorJKHvSX8d7wGwQdJlm
Jo0bQgiP4tnQF8TaUCRpotNm9MVoC+Eg6P3rWgCG3YiS83KpOyKtiUQ3E5PsPlGH
9fVw1BNbGuDPv6tDg7cjpEWWvzA3PMsPelVBlHgi5C4DsN0+xZMXW8WjkHouyee3
5orywpOlRzfC6oTvtOF9Br5OpPqKgYl3OLaSSot7dzeCIlQRauLEUywD4mGJHnqE
PhOJua5mUBAfCSI6/lZ8W0XNajkU/zHAjsyyg3uN9c6ykd7hj9Ae8gfWaYRuz7k+
KyYXYqF6GePf126BwbHQrzcGf0LRldPxkqXubfIOdmF9dYBVW2V7EEHaIi4lI25a
KJaqh+KyIssLMTyZYSkrrvrbBYgAiMTehkkjlgJAIaCTK2V7FiuEMM4lk5j5bCM/
sVpimWq7VLI69DKxW5KZh7oHbR/gp3UeuFiL144CxS0FIWuzOSYPE+Rvrr1DXA87
xeLmCuMuM43DidTFlRebRGhUSzldoCwZEGbJnjDJQnmeHH7aMWtgndZKw3RZ/UTk
CIn1ADrvuST2BHCoycV0Yblg1mcbf21acX8WKvNHohOYDPQYcYRjcpZ5XvBq07SW
W+uAxQuJ15qbkLOu+w5FEp0s0DlcAge2aDuEcRtWsVasYA2/4hBtrugAoWnvp/jz
84Y6fMkBHxJZ2b/ZSg5V1PxI55kn4DLsDx98gWivZvRQjS0FEWw+SU4M/UrRkbmz
cGFeleJ3DIOCoLjJZZQZbGl71mU97fXS5KPeirkZyNk26Lo90AtUyIyXf3rEDXnj
yIAOfZZJl2FgXPVyYz6x/SvbHyT/+lcOEVzIXAU4nzv+rMgmSgZtVwJdEGWZv1ek
+TvL11+roo9hKKHicO9kQn7/II2dmsM8RNdLBCV1a3RIOdsVxHwTh/3B8fPV5nDu
knCWijfNAPYWQph05+yuJ9v4tzhYisA1eywTFSq9LRrfmW9EYwAVOSaBbipSqNqt
PNqoIlY/994DdZFWDSMaDepoWyTnMC62wEejTkkpgM0cF5mWxJWlOU4zTJ/hVkow
5OYXq5c7GJISmbSgysu63mUe7P+j2EIRNPcVfRB0xkgP9FqAXGoVtCdmLwoatXOF
p3x1DnHJH+pnHCjquvsxJA8jmUtr6DKs8/GkagwMp7wmteIa3+edGOrAxdQ8sw7R
/fl+g/S1tI5omsGCroNnXLvX7b6fWzyk1V/zhJOOA0+79VU4Wc6mn5fv40a8KT8T
B6MH/XkR7/STGCYUcOP7MpmUchfyob6y1nFDKui4HOUIEvB+9ZVaUP+nkVHEnIfC
1/ilEpLKEg0iWlkjjEJvOoCsFfk36pNa/FzCUkVteLtqqc9BM87pWpnD2/86wA21
4rbRanWqsVfo6nwDInt7oxI+51jab6vHz2C3swFIu2EORWpN5+NZEyIRy13EqOYd
6mdxhpqmprxmscd16oMPM9JnyHFkwAjT6Kruo+02R3Kxrad6udAdeiZA7VSuK1ej
o7XyBa6WcpvEwppeKKGgAGbcg//A11+s7q6VR8cYOMGuvDpztxvUJZ6mCUPxGHKd
/3VLy7IBG5nY0UBABsGntlHx1ggJ+ekkihr4JQQFq/O7SsVg/lTofov4rtazHrp6
tmV8rpFiRtEKc1+xql1W/K+SLR2F/SwXw9FnGVT2t7+ObgAOtENlwnG2bRcRXx2i
pEU1oi1ZO4/+slgh5OjncCq+OH6kv1jN087zLzU9cMcDNaZiBEGLeEUWeVJ95d5A
oYDHOIY4oNs7JRZ2+whnOooiUpqs+txmo3NQFu3H43UbC23vu9ABOf9/azYcW3yb
qH+DMmWihe38sL6ETKaJtB2jWlR7jiUj3ywU+hAoUy9q9jN9dgl9yV/tLJKKalz3
/k0Ln6pKQ+E+1lGkLtsgs6TtD5yGFOnB1JfjrzsALf1n+9Wjt14CBIDFgZQLMIVy
LHWfrtRTkw3BlS+6VxveZ6E0gcb9aoPnY1Cxb2VEJZ3lLwNkgOsUkLhW4Jh748Cz
VX8byNyheqMyg6TBfvHlRZ6BnhNMngM9RgXxM8kv6kow9iNKYt0P2ouv19NlVwqL
Ruz2xTeFFLMAg5uZLOTAY+CfpnVXm3JnJ58np5t5ZCWfpPOyIgcbGrK0YV3RiiDg
pDDRCIEgJrmepKK3xA2EYTN06T5ShaDQnMHVG6wwacw2edujk2QFkMycLj+eefhc
aLWW6qjgl8Xx/95VTtenNivwDn1W8bK9uhHen4x2NnCDjmfQZB9LI6FF+IuqMyYn
rDBFiRr4qMC82Ix6/CxJjv9g33fiH8RIGzB5Oa/bdBAsjToq1vfXQEE77jmNoPDo
JClpg6u98fFASJJf06IS8grUjie/lWjxm/ovNS6f8hgQ8UkE4PdvxBjSv8EjyRO5
OozSVxJ9ACr4hwG5UMppObTaECIw5amElXtMiymNAOGFVSOkDtfYzw+W8ZDOFdzn
rQM9xmDHIflhTqNss9hmxVQbxh6wQrZtF2HKmAL9Sl9Q+S3ZKPKohAELTciWmIO0
I9n3G2Purc7mbQzbRayJfU/RyeC7K6IhWjEwJStD3Am1RmF7aGMD3vrYLu+B6SZQ
hfOFOVjtmR6PnqsdRo+bB3QvLWlrV1htYdN+p/FNQNmTFVlP0EdOHd56uQ696Uvw
NJUA+xjNP2aPDjmBdssiNyhYQwYbMGFl+MqH2zVC93GpYkQ/kiCMX68gb9gDo1pg
9BdyUtSr1mv1uDFxWRjKPaIxMJ4QEw2S7EMj8XasSgTqLxJOuSICn3omb02OXFRZ
o2eEzK65JY6rMq6xPaWMODr50oC7jcMylzZ6Tc4m8l7Gc/Ey6HbMZXNOobQCDnCv
573VjNPZGZPwMcliXtL6Zbc1VEpzFgGjkrX/kINzxb5h1/BQ3b4y+vje6nMSteeb
oGQwHqW87rJnGPOrMZI8RmG0rd2J+JwRLJMzNly81wdoPnik2iYGQ6IPbF/Hl64J
+LE7wmcjjOCtB/OEDUzEs0CT6EpI6fQKdmHAhFxFJZhDWlRy6EjxU5FkOuuWsWVH
BbkCt0qVXSj0MSffkgEu3zXe4YBq0Cq1lfgKqr2mlVFT9svfTd8bhxe+G/u3Pxvv
1GzWoRDtoK8wjexgc78Fe1bytwqUZWlzERS0JJs0N+FtEE5ZU0uDpY4SOv2O1PP7
dVHh5mYXr9WBLM3mX2yfc1XVE/9s1k8coPsVpAke+qK+o129DuG5I/DZ4j2T6BO1
P/Ps7T26LNxQy2M0P7cC3YLKfBiDGRIpPup+pBTDIt5PzV0XUock1mj9ZiJffZTJ
+GYz6Swn3D3Bqhlr3zldY5haLe9s2uQB61if5jygMX5EtIeOOEvqc6e6Pm03ltfH
IWJycCwBDmfy3l7jyT6sgcP6wpUdujTUjeoSsim8iGiAw8H8tg4k4dkPXTvJfP1w
dBT6zf4a4aQnYbw/sGzpnE34ewpFPv2AuNixuyO4K74dhc/jWtHpvu4nzb3JhJn8
vGIqndDUykWd++hG+TvE8UHI1IF1ow9vV1CX420Eids1hpznmV4uO/iJxlaiVsvV
p8gKK9sRa06WuRfu2vwYQvd0BYndrZ8N/+CKTDNXdzjKkLQD3mrTX1HuH3YM3ZId
gVQZA4TxtkLwDUJCjFSYDMW9TRbPYFgq7WeS6KQsLoTJUHTweN5PRg8NS8/0L9C2
4DjLIEeJq8O/NcphmQMwQB7yF7NhNBBQc6T9tiNXg3sPB83KysNGLRx7G+R2lcrp
wWJRej74ZsYqetWp6viLt9F9xaLCgsYCQLlHcG0OWSeQuRi0IGWWOlXi/5S5kZCn
AdIwggZolZrpw/DmXdrLsqRgTTaVKRmwWzLzM7lS9UikTPqCaxqMDsl5bwCN9slD
Kz6E7r7enS7+kx0k8L3s5zB/vQ6sqhzGb7BIZRFtXNxUiLGMUxfNiwUXL3kbr/oE
e/PSlaSMDUsnxJ/T06RmX650YPVclxUegXFRhmD+4E19+78AUuBHtQYscnZ9u61x
7ax3FVC7CZXv9sDlYvWfjgzPHI4F670gmjkiUQZBi0Yaxd3X0VON+z75gMQxysPd
ii+5MjA3eEBEzcprjKwcGGV/FBOSV232roAKHu8ApnZ8AEoGf6Ixgmgk9i/hOZ84
FlIjUWDwMlq8Cp5ZWSbayoSv7QNruZxEgFS0p0wjA719bU/GYuQ+HnUDtlyqIXli
FuaXQzK0zfFnDGnVheboEc18XVT/lv8MEoIaee+DiN6cL3CnT0YAVpRWXI4M9QLJ
A0AZO7dh34GTFqRDWLczMVkRn2Qgy+4uTiHpC6pv28li9/W83iaKvP2AAVYX8SjT
+fS3H1Uz7D2tdwj6TRuHf1dWiK+s8V8Ire6yJUHAyIE9yP05WrHTccEjaeAgwrTP
5lM67XivWcwv+HoOoPAhsfhgALdXG+pkSR1GNLroe0HYVawjd/QuyGmRPjDCv3Dw
uL+Myu2gCe6hDkkgYvyFr0RRZxsHj7FkIqFdaOCjbQ+ARTLOf5JvBfCSSiZupXFj
GvoIk7EZ90Lwey8Te0WmOgUg/ZOtSf639mxkWU02iuVv9Pi2aqmi4k47eFrJ+ow6
uXKqV736Fu6Q+8hNVn0eQ7EihqNZbjaoEWE4G5k60Ntc08O//J6vYXuQtHbBjxoW
/QEeRxLfVU9573NvgmOtvdfLd8V+C5iobVzKrdDXxnAL2JGna9D5LxAWdxKb22cS
fP9/T/VuCicAdKmNEJu38vnG3xUHTNJIPjLfyACBj81+ETew+IucCtId1YRK+hzx
3ln5g3jKMH4c6AKtMBH+QMNHkdpUzC3aaguJy3F7U52pNDsWc1PFYPTXBpkb5jha
fbVseFMZTrM+rmaJDHVxaatKbj4MuP0QP/ahvwjyxI11kgWHFB8lGdXtssLBdPVw
iqJf2kOpXnaX+1qvQ/0hz9jk0F9CDJKENjk8p58sPsszMeA6Alo5PhGQaJCt/LcU
DTkm1dikQqrRD5Z0OZS3OxONWs9r07e3vcecgGJfJFfpTWFEffYvF2FxFawfCwaw
ZkZDWd3lZPpVuVTYakxkFG/A7XqPtIYYcALx76qDF/bXYwKIJcpHePVAqhSI2CyA
q+qBY8fJCDI9nqn+JPFoVGCacZzghi0Jma8Qeo82GUZkl+ZA92XjTIBlOY4gDqef
dDN3UW/NtTryHcCOaH8uiUs50h422Kh5W/ek6+2KWCOcRIUQ/y9OxAMfPTc4YIN0
pxTWB26MhPug3qFL0MlUI7neZT4FLt1mVgGoUD8Dg83jxVxjVijMXY/vcyLq9mAV
s/7SZYQpzE3vp4bvwv9YlreDtp0QWL3fMqjRHk2Dy5M4fsgtSRlO5sJY7GjPngI3
kymUcgk1GeUxmBWzElCMx5+rptGlmU/LGFKRVcIbx1NQzB9zeKhnobVXBMhp7TyC
OB0XdvwmdyuMO6ScQh8RCamctRqmmg/2ot53KxKTigLmBlf3NJoGLWtoVdGJr6OU
ljCg6WThBFChOLSY2Bw3vfXb8KHMfx0NsanJ1YiFagDEPishJFOjdbUkDGMGuP1u
nQ+ZBr8XsFZYTWaEHscA8ejSjOVwBTuE+xWf2OXGAS8Z8EmaNGCfWfTmzC6KH7Eh
up7hWPjit2itOGekqqCGwrz5faL5Rfq75NHM+Ggi7aGaKuXIJwFpnImiEdXqu49S
lETpxADNNuPmAYlHq4md2SOz1R439s4tPBwSUCrBUqlYu3xWnRoh205mCyDfthkA
SdjQ8+PDUkCy7rHZB1MwTuImM/nQJE3d8d6Lz7CRt+Zx2BVQMc9yIk+6xMq7pL8B
DJkKelG80veg/KySyvb5yzgOGQ0e1SMsyvrgWtVkSn8TZqY05/c260MHtlfm0P2d
dgMcCxfqOVUN26KKyO5CF/xCLJLIQU5qzmAZK4h8e3zAzlznpnzZ1PDtYTF735iA
XGojplzfxL8uhPmhaL3vliNXd3BpO9P24R76oTUf040Q13YxBL4VariCBebx9PPQ
YjKOG210BZhTtzMtc2V+s+GqZK1czFQXXxgC0b7/H17SBbtqSUCVrp7Qxj/cewiK
vbWvSYyVaLVikiWdD/kV9dTQJ+tGOVHeGo4BPD1QbDzTzdE2zTEkdfw3Dx5649jf
q60M9rNZUJPp1btcQj706HYw95j/BCHGlhVR9yrrUTw6OC9h9/ShL8v6fYlM5mP3
fj3q52WsVeiE0E6+na8lxZgHEO/9N0gz4HOK2AqAKoa+Rze63JkfmK1A28jG6gZ4
w7EoY2jU8O38l+Lnt+bH/osokPKa3gJyKtntl1o71Vf2Xy/X/TgvRWYXHzv+20Dp
zqHogQHLPO9DvgjzH5OO1jls1wnfgRRXbgAJno6wY1nWJGvxOVjoRIC+MY7Ft60+
/kbc/quR2qHcGMDKDjYFnloBO14V8An0C5ReQQ4drPCaXvc1rYL9MOEmkOsb0Mkn
6BrRoLJdORhpMWzn7yw0ED+n63hpIw3/mi5Siea+uulDMZWDV/mwTZ2rIM589Xcc
FgDivri5CBTjBMBq6Mml8+U686PtwVKKo2Y7AeN3ADNdp5peWmJEXrz8AeXKb2ca
okIpfZsrNIT4Vhm426vQ3/JrMvurNX65k60WNEdysBV5Fjj5FIK8nODApQE2V6+/
pWaQ42WPoAm2RT5M4stZGqLGNLM9lsFVgm1wSKucixFFhyTilpt8yVYID6uxZjhv
5vjC9nve3bcgCR8ctHgBNqvxsA/puFB0gPIoohoyWm19888ROpBBXYRIV8yh2oR9
uQihBKWjxJAvDpMydeoPWx0ytopswL3duXKU541AtBsP8CuvC9ozLBTQDqFlK2a7
evp0R6ECftcMvH0MWVnOCS1qWQv5p2rprPfEYPcMxpy3sups/ZCchhgqDMJVZw5g
DC8CbEPjHsBG7Mv7kY6unKQhUDdVEeRf6s04+R5Y7glzKOR4jSwVzAWf/IVrF4kn
8o+y1lfIgrCIBUWIy6LqhMb3dx3ab6nARKlgLV5v7yVLNu//w5juF7LKAF6KlLoy
R/yEeteyj0ZlM9v5kXTXgQo8HPsf0rcHOsN2SvHc99oGm6UqMkCa8cVirdM9cWdZ
X4vA1ywuvOEfvcj6sZCM2VaVjza91G25kLeEt5qw6lKgZzxSmiev36NpQe1Cln7R
lrBuFDLLxpN9WwmhIT8OKk+7PZjWGY9UZ0ZlYZiMtwXyY6DMCnjU656v6MS41Q7J
QD99EChdE7dOrs6sKLObYVlWCWV+LbomIt1f0Ow2TQdofVyGTptrmCpsa4BK05tb
3YY/84t5lsfXWvLuzUPQkw/D8+UbrA5eeuKKSKeour8d82FUXaz2EYmKukCLpjfG
x4WnAK12KFfq1GGZc3rlHwsT2bFsNyC/P76FBMW7GbPXw8I+fYEwH8pmwMpqKFVY
/UntLZ41u2CfVlcOCYPxwXB7JgAmWZa8FoMHxAOys8+Q7CJ8Ez+H7jaPCG2vaQ+G
i99PXcYzADkH9qQUiljdB296UziCGyV5v3ARcRnWGkTxEPapa9oyzlhhFTr6tazs
V+lwmx0Wz1GGtLKr+xYgssZBCLkXsXgcAS3lCFDGg4lNmKh/Phafk1jEdhBlqAJl
4G5Gk8ipgKzCeVM3mXzlKt48pzt7pPBkuF5LYIuq2JgiOb3bDRu2bSb0w7EKQHXc
Wk2NCyVmlqef7v2gmtxsp8SeWcGh8apytrV/Zk787SeFrdJcG0b8j5i6hEgIJrWU
wYOth/C3Kftv0l01jmGKKiMSXba4qp9lZfrqxZUYCfcv7HmhAlWDUc0IHfUD6y30
E2n4fHtXkN61R9pdPvuKT732PVrlEjzq7HazQzxfrgD4C4dVzzdqnk6Ax58zS/6X
Go34TX2uRf8n7HD4Ww2uM7eZly266vM5AF1b8W4IHfX07U+tEa9T+sP3oBHLgdS1
fbzTdXol066iz5wWDM/rbJA3IVnH8LWQT8HgHQKYG+RlWUuPNptu0X3H7kgoweSt
YMPMfXXsFWrjrsbD+JeHCkgzbKxWm2nWXt10AipDJiwo3vvSgK2pAF7csYoEY7IK
z/JN9jF/p/1A6QLyXjWSB96Mr+5bFCfVCLVCqoDNljidYHRkNNoK6Kp/KgwSr/9p
EQ7xJdKXlo/jme0DFAaADBJvZqt3bkMnwH8i8SR1f1MD+yj2keZ/3t10DrYEGgHi
ND33x1lyCYFK/RCt3fw2FqLnY8yYAXpG+UxhlJT85O6vESvh2UmA5TFQ1XBlVtju
y8JqZf4rJnZXnMX8iGHPce1/o3GV98jQ5AUPe7OEicqwRn/nVU9YK2CTJ9dXSa21
RhY2hlx9MHgLHHyMTCiEK8UiJseBv+fz3DzIElWgLU8NO4PNrh+VNA7d1gD8S8JQ
IOC8SjhcLPUFAr1AOHVHiJ6M1phRog0YXzvoNdNCyMvseSvw5af0ab3qsy4LsVY0
/fiEJo/CidjUIiTB81xm2WkSVDWEmrdfqO1fgJ65Zf/SNa/B3A26OYb1RTJVEHIb
Eb6QvkUNbsIUyhxw6MICtYXJZk/+drxKspGjU4ZqGnraFEFNwfBLCsg2hgm5m6oZ
yZl+/md7iqsFS/t3MFCbTaiKM968Thnp2VdPaM7GOe/5K8SGEMKNy4d0vxEObdpF
Wsqo9Zzn+7xAu0pXUBXxzxnxvmOBWn2uovpKoTi+jjfkaZKAwUZX25U+TvlD5k7x
INdQySc9UpC2aQiK0qvCy0DsPSGZxmLmgA3MYUnjNTptRkjm6Gay+61u2EkAa2t1
MYaJhCMj7hTkflstsWWaqb/jGimNt6NIDIq94nEi9L63Z2aKsohcXpnu2msOCKVa
vRWR1PEB0rVTiB1MA21WHlbPtdohC5unn69vIODd7Mc2XOXOgAdm9EOazSH30SKZ
nO24dJL6v9TYu0uobSjJ5f/WyencFiF8xFvAttrZCmaVf4PffhJRCkJbNNvaXaX0
pPlW43Gk4SO4rNFWE5/i8M5XWA3SC1Kz357QS9ziXbnchOl/mRlvUl8MpOpiVBkk
3vU+jOC1ULJRBMK91wOi7xLgyc4bpC5Z7LpephtjJkdn0IFvBpODXr0CYQ5McJPQ
3GQiRZrzmqwEQ2QEt63hWT9vdfm3evRbCexkh5CyYKqj91gnYMcpFNRAndPN8K+W
OwryvZ/bUFDZGdzLCH60He+lJ3q6iI7UHC9yRgmtKaVCi4VqqNZ7R/3TP1GRkNYX
qY+1l71fcqiuAVCl+0g2NPxxsHExIBxODXSYFMSdMdauEdCUfupM4Q44isbn1BV/
JrdcvEHV8C+zPF75Xfnxg20iH0leFUVIbTGv4Gr8OiU9wawTDURX5BT4JqX9Xfhk
345MxtOGTHWEIeXYl/Ms7WwCPuppmpU5v3M9nN5EO3HdPvK5qEjvDhoUNJGv5bmu
Ky5gkdk8m43MtTLYPVuNeqc4TVJd05vPkplkjAdTvDj1/MjRvwTlmPRC/WzC0sW8
t8pXxEg1ca2qoCzBsEA01LqnIuovyUS9zuD8JszHDc/2OLHxILr8FriSwsRRDFjQ
5GNJAvQ8ZFWkbOo+MosFvUK8BPxW0V51JNNpGqYp5Oje/GoCcwrkaxhvio3qdTAA
XgdeKmFOBSnsNFqdrT0V7mL4n8cPESgmtQG5B8IxH5PuEq+F9ljhXNTKBE4V7fP5
s21iwrt1boa8WdBiMHssyigdFGH7RXEUN1npOuLvhugMP+8tXM3eBsjO2azmySoO
7HRohfHE7N7xUoP6KR3dhJWby5eu4t0cuiJLsras0avl2LK5CJy+WLr+HdYaKlBy
ev9U8lm/oapicjH4aopFF43yrPtRuFXKAW7rDXhIfnR6c3W0AuRrkb2lQcon8Y0a
QIQwiVQ3cNFiGLLHeECjlRBN4EWQ+yX1E2NhdK1MyAZ8oliZtq/3GIKYegXU1Uy0
4DmSOykbx5suWVRwB96ErstmGSJGSfplLiAtiNUZw9UrqP7LyJK9S6YbDdyD5CpP
+9TX0dCiz1qvdiTUCJ4B+HY3tScjMuGDL+wkuiti1T7o4CKMFYVC9fJpGFaNzJ0N
lavXAicaAf/mxidVWHtGce/FTAtJoae/Lbib8k9hgcUq6wMtn/A9xbmYC11uLDzr
OHyIgBJYMEKL0GlnLbIFIXwL2pKh4CT52IIMafIUj3eMx1ikcp4zplfeLcVBxQMC
Y5pJwtGh2b27xVC7j0xH1xX4HxQ1YU+3ZfT3h0UZVw44FBcii2FHdG5h758tZhg3
6kM6Ka72+poJL8gd/BQabCGV/nYvwFkmLuF+v+fNRGeDo//zbOjSOG+2SRtrMLoR
usrl4eRE756em6ZUSLPjNgtTFTIjjLPxfH1s69A+9v4ppc5PHFMlmXZ0kkbdWPKm
8pLrngJRo9h+6Ezm/3oMQ8suZLRD+rrW9TZ15AZP1Oe8HSnNclBnmT+pSlZFKLK1
x+1O7D5T8kmaH48MTBFYYsbUqnNYobjr6fcvkiOoNvJXVPKnciNFjLiW0ojtUyT8
87l9lcynjzuYf5K7POqzEqOLm+FHtlKYtVsVne0japQ5E2p4v1rBtc1amFC9FIQf
pOLJSSn6NjdVqWnF3AyGINbilC7U/bfTcsSdqXqtEKtvelKxa+h8Zc4903ru+MGQ
l7W/Iu0VJWJq+xQ9pDDvStSSsxfltK7do1ZPFGiWfY5qT7Hu7I113B1UyorqKV6a
GzbFK+2ue5zEtNkicgEnqf7egjTGBO9CS2ChADcbuKAgF1w7o1kYaf/0Sv07ejvD
BWwYpr7pp+t+gDKxpaDctB9/QOUziw0uV97/bcA9UkC0Qm7fnTvXJ1e4fuC3NdBW
x4zdsybeYO7EG71HjZ3NpQGSUfS4jS0Bi1Yd+R0D/QKXWrKVb60DtbRtUxgTkQ+r
vaCETqJV4CfAlOdfCzaUzC/EMvue0o1bnpPnQ42alp7goQSbAu0N8Xk8Vvnm5UUZ
cnDVz8eiGloIhNfvOATno/98KROBplQ1mNCKZxIqpySVHl8itWtGrpilA76sSn2D
t/8EITnEwz7Nna6aq6Qfnv+gBrJjmNXc1rLiVR1qRfNu2kYjq7sYjzCkyJtKQr6K
1u43Qs63vxyND77yUpdSTosjkz5W6swYZsjcbHcDjEHJ5m6aq3FMIs6U5CoMKapJ
syASeRM79gN4FYaQ7vdZ4GNv6ewcL7wPGc8M6fNzUcAgzYUJzH/Z9ift2A3MpE30
wRj4KW8EPMUWlIkWthhg2tObe43UtksozrJBgZdSgA+NZIxF3EOEvpAUI/j+v72S
KFWwK9guVcAxBZwCcwSYtYd/GsX8afNzfRs8AUWfWv1NW98UE3B8wk/xKvSXmVc6
YfQyctGQTI7YGEF/VzSSCu8BFBGTpOiaJlXwF+ls21mxiQUDFbrWYLfoNF1UNEqg
s0y7reiwJc4apDHCX0KhZjztZ7H2laARiXrzMTFvPe3eI275sU+vkde6bcpYsRTD
tRFaIIfZjXyr9nnp2eX3gVzZjqR6uqv7p8NEO9ikyM3UOvMbzyqK428VA7tXCzR0
ZQjh7aURo+dCnMkYanBg9e9ROAgWfUuXRAttgR0G6Tj7LQvK7a6BQD84EJrTRdin
X+w+SHgjMtyM4mUc6A4YxyyBVqt5N2w1qy1av3Lqf2sgp3wCYPiE0HwQkFIYH90F
bcWHiUk02IUQeYjl7X6lzTkvtjV3SmLEEs2Sqmuff5CuK/HQlYtRaB73YkMPBmnt
FIJlVLPs71+N0gPM/zUSqbVxIDXekIDBJNb1A6a4NX4JCPqxdwZAWDfXYUH6v7ZS
EKQstN7w4+TvBYMO1rBiiBFHZLg4bTuwP90vaO71el3ew1FJgXXmXaGsxppk8SYk
ncyaMA/7HqtlZ8Bbw5nwVUSGN2lKWSf5bNN1qXR4xNZaGUBVhLq6174m65KodaT6
iMAGBb5dmNfmhdheF8yyAVLZdgdFpuUyAZKy94N8vgZwISITE2nRR7BSMIulWITO
ZUhXWhTRTbbLIG/S7ho60BS+izc/qm/mdb2Opbl8ukvptmm2VsWkWpDnrRuDEZeg
2gvNQyRiaPDEeHdiaFE+aW3KbYK8hAdCQ1gpoXLh6QVqexueTLIvpstI7HGn02tA
6wAqz3TwIop9cUeYn0RNxRNFyhr46nElY6NaCbP76xOm0Jk4NOYIQf5+mZEpjRWJ
prYmKjCCbyugLqlKWurZKkcXpzB+HRbvFXX79TuRaQJKEMNTBPwvJNWWAKhFeLlZ
U2lNe1UwAtZFbFx4xPM4om9l8bLBBcclaYtpYC5ZtSRmfCGOy5zV/Euh/vCde3U7
sRUKDIGbdPdq6ae1EMftfLWDKP/EUsj0eUMfWvTWDde2B3cGCJxQvLfjbzXnUBWp
hXV4FSLHRB6p8ceYOXxHii38JEwLj1Ukvjpj1In93atBI4be+VeMh9LTT811ksDN
Xottb3oktK74A05ST3PjDpkqm9Nc2+Tm+VBjKyKQf5Gh83jxn1X+muN0VnKhpIXM
QJPGNNqeg+tVUEQxOax+JyxdZ2VGHrFlDMV0R6sLqx7H0tIVGjj5p/iuFY2mvLOf
7z68xgolzU82B0cjOfQG36TMptyJmeTl8yyWntXCYheflUFM5TAov3HKb8nPBDZl
4KPWdKBxqb2qQLk9j0qO2NM0ZlUpNQ1HQWpOx0IjdqyXlKHo7Oi/N6/X98zggpze
7IVw6/yCJjeOzv7+JWeWDkznxZsSwEqpuTjnfb9KQEqYXnvwIatHO06citIT6dLk
yRv6hbRhuLoNgtF87PLZ7SzcdL4/l+8QNGb985sQGGdgwosPqwX7yHIWO/pIw+XR
z9vhq40rYdnoXJPLoEr3D/qGwGZEnHvIIQAfAT/4DTGkZ61Ydy0gc6zavGRWiwjg
UDhn6JY3GsWl++kjiGZed2lntKgy7xebTUAFFkt1VsEjanBewztOSW8P6IVPPHTw
D+5Qmow02H2Hz9RFQ193GJD31yqkhLFAkgQ7QX1RldXvRQpVA34rUW3hKx7/jK07
X52SMKo6TL7WeBxwMwlD+f6yDrrwRfNZ2TtJqf6ALwJkFFW8MVjc+os87fLLLRi9
tHIsAOGvG89iWqkm504/5jWdWyBBhk57ra+VfNeB2qeHycRdhsMOJyOeok7h0Mak
Px30b3/le2t0E0FSRMfgRinWz34geXlms/T93/lHfc6MhZ8v1ZNo7VCONkdXsv7k
EJbRyBjkTQiWqf80RSkojNyyw7uf74Pc6FhsCXVSi8Y/+o6bf7PFKSZRPMe72LYT
X9O1WpfMN+bsjiIq1wTwdjgl8m5tZb78LG7mjzB6wFVRN0cH20TKj47S4Ls/f2or
2JRtgBSIHiXm0V6DT7ZiNS4Nl6fJR3TbhUHmTz/1NLBFj3ld6lZ38V6gFAOBrvCn
F5hKWlr04bSOxQQ3EbhjO5xtaK1mJ79iZLzDMoIsCUEyjg4/sLHroEUxfCm7hkvU
9VsUo5PGB+l8tp+uugI8/RxT8W+o7M1OHb9ybXO3qTVvgzGeTK5rJEcwYgYJYjnU
Ym5dkxT0n8wLuyxFp2o/05AGwHufTESe5l3aQiZHQ/2+CX6AqoUPQ0GjZCNBYM34
ZSHfLVoTrezS2FhZHckYO1AdQW8ALJgcwxgamrsXZWSyius7ABUlovoJHpKogkOk
f6ZvBCV+a4cjqGhGgv2Dtj3Br1xeHnX0NLADMCJMCn0h06UAAmyV3iOmJUIyRLcY
Ly4NXDul0yjtl80XIcNjA8tYCppuFUGy1pb2jfoscDLm1wFObB68U9JWL8i46CcG
UIK3SrobEeZilPYpgRz6JrbMy4RTZw6wHBeDlnC1hHIb/9yvE7MXqr69GIBOucr5
l19imkI9FzmKMTGL2zFJIJAogH+kWPFk553f6xbi+6oy4pgIfYcxn6/SxDF16ru/
yCuzohaaA7cnCnUuVJ3JOsZDcbRe63KPjCoDTGLFeF4aJOMcYysj/TL4AocGTQnB
/CXJsOx5QcBAXul4ejTBjYZKuhpE5ElrqgqNqJSAXRB17dI7r/x6dG/SUKmrIogy
OCgbgcHhdWaIej9KSEcf12TKgudJiQPtwGT13x3WfFuUY7HfnOo7O6w3EXtPrUa8
5rVT6EeB38cavgwZvUwcIwi1nvHryBliPVmJmN6Yu3qp6Ts9db4bg0DzJF1qfUWs
LjoDOjjLPCPPBDinmKkvlPMbrgYgF9T6sOK9KsaFSSt2JTwyTgNi8W6hpRRR9gXL
Any0H2/1Q+xzqehRQbOKdmLLGAidaDrb2+DaQAqOStb4RL+Bno1ir1yDTjWed8hh
B4vJ1VMnRvz7Ds7m6nZBRXbJxViU5i58tdMDZBuSOJ+YROkqLNFTxrp5Sc5wGlCS
KS+KCVPIGaG8m+etCt4i6J7HAYNY2udb//mrMYWCkMqObNRnJ5s2B8L46o1sdXXc
ipfI8c73Hrv3N47ab+x3oPr92z/cY8t5YKFMqe2mXj4++R0csntvPDd+pPzeCqm5
/i3bXC8I/R+0YxWPCc8AsvK3KFRtTVySNaacBqJBO7j9eW4DXlr/n9tmVyzs8GJI
uhFzDFplJp8A9/daptYAn8DB4J7WpKFi6ngcp/IrImjGI9HDMpCqfvRf89j2yrI1
+ivE0Fw6ARO5AOG5CjLHlJ1AdSoD8wfVB+S+DAPnarAo13hJwdZZWgdsuCo2t6u9
ek4UgO5uKmiyunPlexFNZl2gF2yhNLKJtlbLWsnB07Gmgqeec5iCT/1VzDAKDD6A
rbPF9lcqlCvKbv8ZvGI+p/NyfGZCrUAmYnYdOny5tqlHodoui13LlLOCVk9UJl5k
tYhppeLnSiAah4xhpxzFPJT0+75qrEuC/vX9lWGveI3tTeNVdjDb5eP10aKTXmck
C/AqjuNkS6gluwQUffCObqG12U/JqkyXyhXkP+zWdMRN7Z1oAeNGnUKSuTKI1qeg
KpI84nb1Ma1nk5ZysbHJNyzLGWwo3dngUup1ttPwZI2Eo6wTkVSSGA1qxdrxOfgF
jyPg0Ihj5//Zfrw0swuT0Vm6XbAc20cHqPjamYMlwXUBKuNGYjkkvhWf6urp3/T7
T6ySfuAORPTZm7msnN+Whdh+IV4rCYKJ/k8ZRrMrp6uKlkQD2cK05r8qk8KnDjLh
PwRBvSHTGrFPfMXD+Fpgj5Jk+iIDba1ty4DC9Q+rMZSRTIenu9/JKZ1BqcnOUwiY
/zI0+3NUPssCV4erVP5UBojU8DNWRM7wEXV6/+Wd+9tuE3Sh6iWkRRVhD8oCgOrU
SMLmbz5YkOMfp4PYQvJKKLlHvBnMowTIA9glkscK/luk4hT34RXpRk9DvAtmI8r6
qDqZtSi5KwNYIPv7nQu9SqgEfa2gGTsbms51kv8iJBgNTdnGaz7r1wmcVruFpmTK
ShIQZp+TrXeRaTJuwqPU/mlqAo0BI9GkOZo2XvrElOrvu7t+4smKUpQcfXEzf8OA
EChGcfxv2zg39pTetGG1KQglG0BBD/NsNSMrDm9Pq7rfUJRkMgl38sHt9eNks+r0
f452XFyxWoO3JFCUNprQPLRjDUROHF9lTNiJxwlRbBzTeFJOEAfdTlJtsU6U4SQr
6tFqeojTOeY64nz+M2VDGCTOd6MuIGZ689Y3AfpOx4ZcrDh/yRKh0Ri57JiRF4Na
wgZ2/a93soKgJqyfIhv2dnmr7nfHyT75szkZ8HBguiDxGHkCUj6x0ybUY6r4/goO
3FT/pLw0MIPnHRvmXQyWQ6KXoZkSfAEuM+kxR/IZr28B2Skb9AeqeGaGMlNILTC6
lGXoYyCsDkgX9+SL/ROFrRK/kcUxlsV7Yg5FkIMIVIooHihczrtlpFVwogFnT5Hd
EJWWNbc558RabYiI8googzGI03IIKA8MMXBocqMJz6jrPaEh8KQiXE2Xsi+82/Wp
DV7njLh+blIRbpZ785Ci6PzB5wZGNRH/JgJ1nibyH3qTY/6yA21RMrDEnoNP2b6t
PQom3mP5GrGQod7+RxNXMbqyEaIcMdoYzWjLVtPwpaIjg0kiIZQ7zft8sKthKVvH
yvyK8uc7v670LQ+VzZqhGxccvrH1ZDfta13Y1SrSuVQmnSzSp024+zAyUzZA8u/U
AdPadULRDckA453e8HCEQUEjZXh/Bf95imYQAD92gomkmUGJ8TLqq/fEA7Rtmd+8
mbxGB4sTp/3Asi4RDNqthmZsgQMgnAgkP7WyLFUS+R/alMYw2NUwFhm/Wv5R3nmc
T/PvT1pzDVr6JV0Le2qyeRrVjsEfll43L+YF2cyxWrknihFuVwfoYk3IxDBz9X7x
52CMzdnsj5a3kn7ScRE6x7eB/ow8iyia/Tbz2yq+M96fthENRCP2WIuf4QDtdKIb
15o9z0ZWYbmWsYz4hbIiiKrpb3BRHZPniBiHWwdRxoIB7Z9aE5DEbtMl0VEEcqvM
6fq1Z8r18Evvof9HR51LyvcHfCCeNi5I7khVQMLCEH6/KwytPCHqEDD6SIICAsQ+
Q6ZlaDPssQOBBtIvrk8Tof7JT7uUQiByaifKUawMasXgy4S3UC8WWC8B7dJc8j5H
uR10RgsQ+LW34WvwvK6pNKoYJi0CPDn8Y8Py7+Dt6KvYXFSU2GrivJgoDlv6bVRm
EA8xHYOHa8ExVJkXXGo8AmZm6TgjKNc27EiPYffIDcxJ/MHIU5JhdqLjHW3UwqgG
Pe3ssOJBn5P7Gro0uGaGEita9Wi6hJhFRbHgj5KMq/DeIjYYs6fc4WKDP/rFXXvX
d9bSDuZO8VTTUlaa7s2RR19ht3A+AgEDBCHfz+iE3uyIjRSf82sa+y9sh69tsHQm
eCtNgsFgAtk0XUdXWmlBXCQeCrrAHg1GuXz7MmhUC+yhiQEkrtrTe+cbFEIaHejv
WJPyAe7romZwH8sIrew/FIuQ+GI1nEwqiIu2l/UeFmcuvS1l6WeVzk3afMpOU/h8
bIPasXlvt+ex/GFblyEtI+MqLMFN2TOCLAeC3HuOmJBa6N7f6t56Cm1C8+PIPVx9
R3HZgESz79VGOOXe9T1W8aL6pTyW8sgthLr7XjCT59HB5xVAF7xpf0JO6df9ynFx
XrRO6b+39z5Cy79CJpcebWWdLZUIHzTl6NCyclfZE4r8ZO+DQhSL/aFd+9scD+of
KcTPNwBZnIWCgNvvrcaFM38cXdwZFuBEEOhstFu0B+QchUX0YC+Vypnp7rVEGFBH
cC7B+sGsPrK534JE2+mjlTiOS1DVROuEzMeHG5khTr4sN7UBDSfNYqmyfrJ7nuLL
P+1t6Ra+9uqAOv9nANSzYOyhteLVj6mhLLyt7uBZe8uw/hx7rCwZvd1uPsQ61ppM
yc6Xfinfxb5tXbgJsgIZHUkHZI0/6bKnU0RjXdOkj5tB46ASCm7xxMxDXUj7mdMC
hKM8whoy3QfoEPg/PyU+U459/n5VTUCPVc8EXfgGSJeW0AJZrhWYbyIXbAszCbTC
2H3qMjp0ourpDbzDO7kMNSOf7BAE9WXsJ2W7jorl9MTLgHyjF1rt8/W+z3++bXRk
Wfo0+Y13d4k08flEp3oXOSZZ3TXdRmXqn8DKV1CgUfWXify0iCdAag0t07F5Mx03
VEITurYAQYnwJnGbHx+135uualuwSBSdDEeoFIpQmh0bou/E7/JaGfKbx5CNBSgO
gvFnZwO0NpIYu1Gv5tfRpJa+OAi8T4WqjcgMlXzaIkGndMz/jHEblAB26XcHANGR
e4qV6oBYFMS0IMVGJYbN1fNaneSHhMBLxE+sj4cXDQl634kq8jbRU750vHMtlVu3
hTtIkxgrxDp2gcJxDDIvvUmoWlSbpM5Ct5R5gc6412gNF5BkFZARQ4QKpDT/w9TO
7NfLo3ovs49tXruwTuLwBITy/prrUmXGqxjzfpZ5HJVrhO1NBGNnVy+co0xHjsmt
iKdb6GC/l1X0wrFJvf3OvucpWDGEN/AaQUPkjQg+c34HAtsJAjw6tqu4obG6T1lV
llEHdR1xqXQFJzOR7H/1Rx61Dd504mTqLr5Wd19sAMbz6BXj5FR+bLrz717MIEYO
+MH+84IQXBQFlVXZNVkn/pbgV5T69hSzj+bbQYgdI01C/YWsGsW/M0nhRYtuvnH0
6k8YjIRfSx9qogTY6GYeh5oLhePAF64BDnv1Gxo8/VGKo+AIsNB6Ai/EcZKIediJ
GGvucbEI3G9n8HofQAkriIC6BGw82vwzbkRvK/0VOljRke65QwZSBnQpEcJQnfXL
wFjk6OU4kiOjIncBq05murpO4poHoBz2g+MtC53e/n9kdJ0YsBqJHgpJOmZhRrhq
B4Pxabn6tW1VcNqnJL7hX5tIizbCKKxl+eV0ar2gBNMVw702XHL3Gvc40vrtFDN5
ZAoAJXe29tOW/vMg8kzIqLx4qTB3TCVDCn6rMOZLj+Gb6jYJTMoV7PzYw98rHVPZ
PTCjh+34V7esrIxeGMS5wLaJm57U+taTymjZeZq8tfGLS44VUS5LfTCEhWzOkQGl
mA7hMFAAdFIw8HSzRNcXx2J0I8P7HjUqFj0PObXqB9NJ++h60Z3j46ZK/oqhFyjh
nySERmAXk/zQYsiRkNUj6cbVSTbe0viWwfL93U2XlgE+0numCTurDt4RhyP4RhKO
1gzGpdBhs6f8RU7G58VTBNjIXY90164RTag2fq+h4wWGmPETt/o1H2pPcg88RYfu
S30Li0/nv694aeFmWIj57FTa7GjlI7s7a9f4xPbmB2D4AK3MlGE7spZL39VLoBu3
KJJfazGsUSiAHFagMsDtgDUsKhCPZn5XAvcnBtH9fCdocS3TRvflaLBA7UXZStWk
ux4ehIICQZaymgDZ6WEaAQ5lc8vn5S56gdrPwjG5thZc4+jfspmBi7EME+1Den6e
IxqdWOp/4/dF04+gSr09lWMoh6fY4EIcc/BvK370+MirSHD4tigqanpxnn6/h6pC
ZvmnM/KHfgbWwR3dSOvernY0DZNASXzZWWNJxc9AoTEH1kZ0l832KomUgWNh7iL0
aC6pBjlZwo7Kl7ikdiKgGDxbHOiRFRd2ho8q9nUIOCuxSdDZq8Wn+qutRXJBe4MA
UYeQG5oK4N3Rx6MYHnaDAiDfk/CJkuO9kFBvFw/LDvPGSs5YuG56aWZYEQO3jI1w
P6g3rLvOKYVZD00AU4vX+AfT5Bd+mQE9+8V8zfx7gBS2OZfQ80Dkh3xhqE0/O4Om
ok/nOXyh6oTQG9RmK0vE7X9qcO43c5PKmhhPM++T3Ojg+aygbZYAD8kS08e7yYta
G9iW2IiO33VdY52sFhTghY95dyulKxllhBcfoWePsn558Ym/TH4uSghQ57chckgM
EyKdwIYosbG1G7LZpysm+UleR4yb0o+9qTnY+A1ZwqD3ZU1klU5Lo6eBVSjnIAwC
fHXNPmUk2qo4Day2asEV47uFsZLFa2xXYeh/EAFyAsadi/JeYQ9LNcr5e9lXLkCA
WkqsR9C63KsHFV1wz7QQq9fJYh8Vla0SwNceuIovgf8GHl200bu7fgd0SvMIsxPH
eidraYWXOa2xIOc0cnfU+7XIvJCEBWhb0VwxmVdzIkPjwfE8yuEktnJo/HzfarvK
hp1yEmEwzYGxlY8JL0Pp7fkQSEPrm0acYxmBWZhciPvzzRScSNEGArvfv+yVH+ue
hSyZssj8RjTTFEOyVJZIO2k+LOFKT0vMpGcaVuuOoBxoZ2tnBb3rtSqvZaoeUFtJ
pTj1gVGahFQG6amjVwogGRd+cDd8guIrxdhvEkD2I9MqvDrHiguSGKyniBLb8x0R
l3A2ZP6m8OAtaQiq8JQvldcSXKK7feyLPznRm0dKjQ1gsO5gmRNjeLiVvaW2PsfV
M5RHJnSfRyTCGQxW0+6tqQIomrFnoIlmK44gnjKmzeWYAp6EVuOFJHUJvBgx05bg
drqHqinaM232ey2WsrtSnAcxTZQnImO0JATDMB+tbOVo7XVPpHyYgjHv7ewzqW4n
nH3Z0D7MvdUbAanSny+Bzve6DFOOjZnHiOq9nBsI0rusgwZ9LVRhe3abbTuBjTN2
U+2bN28emFQPrMi5YBjLnbPbhlgHWbEKzvJGluNTNfLEBi+2lYNjkowss0zVTS3x
fG3+tt2TJmfx39+1YvW2PtYMPZ4uSimYl1JwSHL9vvjXFF9E46U8Nh5wX3zqGLAQ
prsLZmtM/LFLTOvaeG94ODs8fDHNIFS8rllIgdl1UGnmuskTxqpo5xNOueTEOJlF
Q8uvkooR4EqpYw7YVPP8GUfUTyLiuCVXLzVkszW8v0Z3GBI6B6imCVTsWYFfbY2l
8Nl0xr2aYFKXs6q72XBXi6Ov2jFzHaOS2UNFgtoKJ9g4cmj+h+uMCe0zveaBRh5i
HrqWIW/NAAOftBRk7y1vw0mRZci+ooX4RyvDwCkUOTX8wvEW3qhYtc5z4j2D7vaq
SdwRhkY+caxD9C6y8B8Y1lKSxgyoKKvWRVYNdE/6LOAVAGTDUnoAlMpMFS+uBzFt
V45lzjucU3xEB2O7Kh1pC2hwQik7dNF6lzPtpnrRMnhfoRKcIk1wsPGTT7JUaJBf
q/XZzqwrOE58ErIA1HdrwSgH4Gg7hfNTHNQpMju/t+SMk1esQSyKJklRZd7eRQMA
McoYlPYFr8hPgE606McnS6URBghIXBq9eTDzZQxfLBAG/8OQ20Q0fGxlOzYMXjA1
zKe2UP0NX3kXKeYptx0vrI2IQ7mcAkgeJ3rlGR2kpTkSLNSX0JBUaE8SbX/UQ34+
zcz0GUTboil+hsqgTuLSPAi4/hsW5l72hnizSLBOaAXqrCNkMvx0wnimRzH8X4ST
Vd4xadXybvDn9UTWrd4T5svFur5LDcCkVPgBx7XkR4ngWBw/maakG/DgR85wYsNg
tSNDlIuirLbTMR/2lIUsnzK0wnPhYeu1PDr0cQkfHH/Hjq5Wo0+SXyeRcnH7K7SR
9vt70Ib+U+lD+e6nwzajYRWLtjGC/2GhRuOhZhyxYC2kuIZB0qWW5yYRrC/s3uCz
X/hT/vvlFN+NNl9oT5lkkzfZHGnKqY2rf3O4hsTDhos4WFcKO3SGh/V7LqkC3bcY
nn7CYRY3J5RTgz0PvmmX38wJ9eYlZKceBvJoyU6sC/eED2i1ov9Zmg8nMqVR1vGZ
AYyWTd3zMqVSqtDGLrANrRQfuI8XwiyWBbWYuvdnw7XeZsZnVSLRnncZ9YeO1vpp
VRjjv5GMlULwUsX5nF3G46ATCqD3EfsFOK8SpLynVrjSqgMPmCapuxvleJpnHHuW
sJMyiUBHdZOWJtY5tc+trK1VZ0M7rB4YRDIbfS/cLjGXL8eUd9kKNfcsd6sd9W+m
yPJMjxTVYD/z5FpQe/DnXdAg/aSCaOjdQ4BJwQ+xMPFGQgXqDHS4EpzkEjTzkaCL
mdBLukmGPqIoCobg/UBuWNRXINH1h/z/DDzaPUa6d2mKM0x03DFVNzSQbasoxvtX
+kCIHodF4uGGx1TlyC7Il5dTlBDhlAYBDhAWCbtLbR2Wp02OMI2U7d1pNIJ2fRze
GV2zsiBUT0QYJqQaiOIrdFb9j+NRaFKuYkSu1I7QnaNbVVwgyzOEkXG1lY8y1zQv
qrnmZr84VCX2hiWZdmF9E4xR5dq9IBYN5jfn9ojvmJPHlwIkhV7iqTs4y4ed+9Yu
rt74EiwlF9tjpD9VdfYFBTWs2/A8qca0d3ZNacXbJ2k9rwdEv1qmyCSfrY4o1CiM
W3ExMKQ/yXGEIM/hJfwiJ4Uj2GtClFlEXpg9YYojR9wAvQxCpuVCadLqpBbHhFkS
k39+LGhZLFhmFThBi/gLuvQp0FWmhHFyfARtQc66hst5waSSQ+85bOfpESYl0n8i
PuPoqFWkZ22le2Ua+9Cvjf30Vz413hYlQxpl6awg9VtLwT73XTIt7M42WsKupgZf
HXlRDl0F7N85Maw7THOpQAEnX/YbiLfWXxDIQpHkJlkLRXP52BFfakxLR13859Pj
ix0J00hCosww2zTGpTk9129LytY3Ro1xHeco8MNhEf4JGlmO2U16098VLFVtxAs1
lWAASFmBaEsQO3lFWcUdgqfQjjKpLbp2J748cMy5N37jSkDsjhBa5NApBtEDV5Vv
xdsEfz00ByayGi31kiEGZ77c/+miKysLFcvBnZCZr5DO40bykrzcfUwl/nLFkTxj
zlWlbJ9y18ZoVmBBv+d+wOVHB2aLEO8J0csBWeuQjlpiuqOYbTnTA1Y7J2WpKT/f
aqhuor0H0Pf4hQ1ntqd+ylE1eZ4xbeI93HBr9RLhhh9pQry8OVeQtThJNw49jUHq
8rFR5lCUkT+56CQ0quE4Yz9eSHl8U4e6044r1dp7yX8N2417C9ccQoYpnuedxz2M
zOaTwKqBoANiNlWdgUqi4NlSDdzxRldlSPSc3kW9ljsRvjcXCDxArel2IxXAVGW/
3NouXgnMdQxkCZPs3hTsQJjhpjfUrkLiQOUKSGzJkb3GQENueM80WtDoXy/ukoN5
jOYgXgxBazM8K6uIh6MFoLVsi2UMxiAogaXa0A63Wzx5Pa0fgpUfnfxzveohPX0b
PWoyYFAwt1yThHAXdf1dZ7gYuogjyTNU6IupRIj49/mTu/kXQkDI8dAZ5M6ckx2F
tXw2O1SZZXViIp0C1rtZLNOHkl6NdQoH3mzyGP3nJm82zS+FnlLJslY6uRhIuDYY
KItTPx3R7AzhCkPpxkb/V5qCET5MYppOwkH7ClOxx2nL1R2ezjId+PgCiZpv8HxM
wOUglzUKZcLdV/tl9FLRUA+bl0OoK8bhd7LT/uVUWsI8+d6b0r1Z501TGz3eOqNn
RyxEfsUrxR+mi3Wflq6w1CsbA8P3Zyp8R2dMEvfiZavuDW4kxHEs2NFLsFW8lya7
984muQtGd+jM5t/uIEnT80TQ7cTGcatjkAfE80eC9w/t/6x/MVgOfc8QnA7vFmDN
uFHyXMIe3UFYZ3mRuDhPe6XIFFq+OjumibYXqBKr3n/Wa2Gq3ETgkw2VBrOXCDtG
V7oDYF/1M9bWopSocrFS6b/J4gLRHqd0jNPKvaTpXTl2us+daWABsEU7sxVJyGOw
fQ7MHp4lNMOa4BpWGT6oMp+SrMU3GV7KlET6H0LWsJTaygSzmGWy3NCPi/ujn/l/
4tr8EVCSkOVuJlbj66t6nu8QTQXr4R0Ne79NppWaHP1gl9pB2vKilXzfUAn+C3Cg
Lud6s8xjuhic43AEYuzN75dXeeeaOkeanO1i4DBYWksj2dBGfPXH/Cahp0Mn8tgi
8aHFoBBAbSw/WGCVqP4vAwVATKkNvn1SIPh4eQmr2LKAB08G9gUNZxFwF++BvIhB
KOf/AkInh7Mz7peqA0tVpYmaYOYSpSGYFNL9RappSyTNMzgBYOEbAjS0GmkZX8tx
nZBpT5ymzukMCDORo1dLHvJ8c0BLXHS1kZXkzIdcYfhqAQF9aQ9OOW5RjpbViDGh
vlCOWbKk75qo5ii37rhBtJtHcy+iqkqJMvjZh2b9kglbHitPLUWlQZmwCmPsDVGX
Y7If6tKVT+J0JoAENDw0OpulS+Fh6Ihsolgj7g7EUh92R+xjRoFhiXnZyrbDAgtr
AReuIa1TqqjbzaUfWSJ5X1X4+1S32ADri3x/TcSmc6UooWziYrHlgo4dzJYUmY12
zHdTercXliy0SfD8gKtINrlk69jpboXJuPQzQJX1mFhaF8wsgC7Ks5XWocT1i4Zv
X5lAfpHDtN/lV3+E8Vz7I44MhPaAiE9wra8DQvZp9ypsVsJ2XliX3GbjUXp1FttI
XURU0Z8dYpd3fjzNdgmrmDgMnQbn0G569eoocGzG2kEItPOHRb7gFrlU014yh3gG
uqsUiahlY6hT8tbVZiz9xjdtFgRthsN3RssVcQVuX7d5+3hWC50v0odWsAiPOyNY
LVms5A2ESfrI92UhZyeT1haF8uraTeeGGDFohCHfLC7B3+UB2VEmHn01RL1hWCpD
mu5NXtZz4MOVxXZ3PabmnBYZpIN2IxLNv7GXP2PP87Qq1UPjgWrAdHJeJGw42/Mv
MitJTU32y4aSW5blcf00FxE0n6gog5mkF+Rl6gQGXtNxsxTwcOEs0O8qZOH8kxMQ
pyvL9wps8ovADfHiSELOPW3wUuunoXuFbZYfOKpXnZjqEiW9Bsr9cqtUIExxsLe5
AZBdaFki6Nh0o2TcFDr+mU6/YKYNdwfwwKee2IeX2scqX3PkUBG0uz5PQfHkmU4i
82ano2NpIA/SjO4umvN+BqMmYW4nDmH4h+RTT+f5mv0LCPrgHkgoaYuIypqf1X7e
XWsXnRlZ+rvLMlVnsuh9/GT0Q8MyFcD0bSlbya65s05HFksJ1HTX2kN7q5JQRPKs
C33CJ7g08xeFkbgfMit0QsuJSQp1Y4AD0YTqW5lq6VURWEszsO77i6sL4I7fyy81
827ZZKQj9xnVAEjdcVJ6X+UCAXDWd/xc0h8Bn58Ak3i8XJm3mO+UuSx4evgO9VLZ
O5uF3xOqdVjJvpgZzKIXw+p8hMS/qyerulmroEqIKOMt+DV9AX5PuRwTUXZHPBDN
gaZu/8Y1OJRGuW0e7Ck7h/jW7UePKWMxi4rpA+KGutvDPiKMHhZ54PwxAd73bSHg
sk+hAgTY9rlcbSczdxYqPYvWv5hYXS44vZlYAi+40VDk1oWgSn9ipzrUTvJiI8ll
48f+1zhGRG0tily+fl7MLyuKSyHxF9qxcnXHWDas0yKhBdtYpLvbyyJl5Kh/9xUe
gAoVoW+1Lz8fk0REy1TWSGdtsUFYB9rprTGIIXFzIDHoriDER2QH4o0njqL9jSNf
D2S3EbjcTShCn2y0X49vRs70k2RQoim7FGBVwvtSIfJe1HBdGp3Tj51gy6o/fLvn
wZDNB2bQJKu2gI6cx1ViyX7YKybLs1GQSKV5fZ2S+DJf4fDa3WmZlgvSOlwwcoKf
U7xm7wbiLadECiGUMcYgqe/+Z07laaeSqwWRrxGKbktdty237Fv+IOlqydWzH2ZK
9BiWxHai4wb9r0pCe7rKpjtGDYdIjhk9OAjGPTyl6qvmxbA7StDT725wz95hMEEx
qariQQljzqaE90KqG1jx+UnfqwcP8AHcQ4lp8hEjVIo2NxjJJuDmtWhP55t1gj5x
DEWv7qYVQl0lM1On1CorbEwVMbhaCkfB6vjBELr6OKGZqMMUTTtYleq/Q/rsT3a1
41LuaZ+iL4x5Jib9bVilRqTKulYpcde84O3cxxdcqOTPBNiEQOJFUyaLEed67xsN
H8tblOnqeAm4W2uY+c/qUX3nOwOQj/Qfpl5Sf/LDDwuMwvCT05iaLWIfGtyImsj8
fl8MIBLcRUlvylvgFanqC9ZYGA1zSJe2o5vrEFTar/j79sK8frv7QEA/A+f0Q+8T
FmCkvGDCFVaOmccg8Ugt45oihMQDF2dknP7NBII9dWOtJJ3tDDLl6zSqoLfqDvEe
1HllRT19W+CFOR39XmOCnisPV09p38fmyV8FMIVQCqw+kFbBWiYyMxsniDjmbikb
fBkn68smQcwXBKcRxa4EhwDJBcokTzv4jaO4kegXE4dGiEQKXfwh6YpccnXLSHbK
MbrOPjWOBP/bIPrcrE7/3m3dvEXCc3SCiTv6OWBmHtGlvUsyj2e7i0Ikw+iMbsyM
GF2Dh5M3RuFjJJhP3WAbKO5ul376zETaPEFDSI7r+nCh1QacoS4uhCKyHzpHy3rE
Uo3NZToe1a1EfI0hbtLxfdO0+VTEWVla1dy8TTuhdo6CKPhOvJWsS5VPqVIcWXKZ
9JTtLlWOD0uhW3m9toDmnYc14KEZZU4a1uZnxszSLV4znYiVjNMIXYd7PgD2i2qD
Rqdc83XlVj69G44/HOt502/Us7b1OsX2WgPX7Evwad76Dz+2RPmC7OzwlK7C8pax
FeuotQ747cswQGmuQjPsgfH4KsJ4+Mega1bgL2klX4DizQq8cPoXz0UUdVrx0mLQ
Wtn8cxQ/DSgUvtr4UvRsvwSkdXAT4gaVu+sbTa6MZnXVeSvwQto5VB4vRurueWdB
3OBJ/ydjaQNd0LHtyTK/MkoHITvDBdROwPvVP4MRZEnlSes3koeJ8B7cAemnNeEG
Nu2d0OgessE9fnJ00XFrWG5pS9hENORgIRS+jbwyAKhy+8wX4zu7Y5qvP2yywIlg
QwrrUI5doDBAB2A8muv4EXr1CboDA44mToF/Hpgj5apIphz+wug96UvtjMeNFLM2
3tFOpaq3uw0t0v2gEfW7BmuL3g891beqb0qquMSDj7eB5sQNLPT09ABc7N4EuxdU
1OdCuMuwXlTgMdrAn0VY8ptlT5OmekzMrmTdJZvg0vfjOdkS0/HNjtCWXAqMmY9+
50hzvjAx0RlLoZQtXr7h/FEzwqsCsjRZbx7O/8Lj9VP1GCQaSTmwlgSx6zopOwLg
d8041ksU8ek5EVpmLNdWtpXUnR0BsqSQYcM23b6U5z3pEvKtcdWzt778Tafy3Max
OXNsTh1DfcSXfUEeS7ahiIjs2CmlTfSOXNuZGGmjHdaqg+ZhaFSoOjXd1WCGdr9J
BfSyo5gwfJC+OPxW8i43LNshpnKjxhxHbCikMbI93Tnw8Pvjuzaznky5l6u6d1e6
n/PkolIFYPdlBzwdjt3yGnkDC7bLbPG9NV10Uurb/EIHRQTynw3HrdXm5SeFLu86
5pfOvMIVoHFZzV41VXAJW3kdsAOgKry5nXWrOIPKyFE4et8Ul3AJuPGWoACQ2MC0
DHKLtqY1zmctnKc20CgvoYJoQm43IE5D/14p+LMYFG/mQ8xj5hMtY1oLGWrHV/Tf
T0DMh6zFZ4kWrLQXs+S9KbS2Kv7uM2NbiXI3w/c3pAP1iy48/zCPvLX8GfSeSkuO
Ie8sZSXSX+Vo1O/eOh6rg4m95N1R3+LpXGhpfwYeaaVIC9dAdu8vtaux9hrz21C6
B9cY+B64M0nEj1F1KYnGYstEwsAZHqUE0YLGk6EwhRlaMnatWBPFX4X7Y6ztVw0U
MipsbFxdtjhqhUyUSsgvKAaYdQKL+9DaoE9u9BY+g5oU7g+Tg76G3hne7qMIacrw
EI22RvDkLlDONFh872wPg3GjGC5nmQO1EebioQ21IcxdVMKNWmBx155pAW2vZq2s
PYOU/r/XTI6trSm4LeWOGMVhCRFDxYGFR4OGqHYBzxIaCMvwbNsb8h8oltd0jafv
p6L3mtaHGG4XD8s34iNWS6h9kxD00crDs/w2BdI1rsQ/foYUgQA9II/hs1atxA20
22l4PHPs5rFaxFg5oI9SyOaBzoJftMfAJCs9xP9GGNEkDAbZj2J6Ru+yftWyoDSF
IF4m/Oc137x+lZrd5Gk6YthWoQMuMrdW4tOJ2n0eMQcjO7JxfgtEXPt6y8qPT00c
hGJP4QiHb1CUwO3u5YV4BWbb2M7Kd11iYVG1Ft7YA2RF3Qn5ryR55Zfxkacx0nAF
pVs4GXPwbwicvoTPz59E3ehfcx07DZCcZocdOI5J+Me54L/wnKGOsvLm6lA17NYg
PClRW6SbnrEhDgSlTZyFmXeL9mQh3uAcJclrWjT4dAQDL9IehFHjrQuCKbMritQr
U3BPWlci2yzHX1JZQ7vTBMzG8lB9AlWfD3Gvq31UT30DLJ0C8n+YD3L/p5cJ92OL
QwOx+4xwQP8350t+nBXrwIbmnsWcGh/Dk5eMMdnmN5pYMP7ewLHKNNjjzuKgjv+1
7I+Z9Myx5VFr9zd43em4HrwhN8qqyEv4mfua4Lsc5GOsqKz9V/cx26E0xcrZ8kcS
I/FGi6NoiH59iEcFVQqQeM+7156IGaepAAQWlg/EuMv9Px+NbLx9RNzhvKNZn1OW
UxiBiMRiBhWnvYdH9ib3cbpEnu+iO/vU08ZSWWyxXiSczysMqLTdGgviQoo4IzHD
1pOL2uoJxbyNkJfWz67TOdG/Om3GYEBZG3bUnoDs2yHzMrBF8ZpAtP0jIIF8hFQW
/TN/YGWnclLa8PXH4PPMAhp2m+RAgC+wWwr5di6ZkfMVAa7N4wZ2XiEupD3ag1oK
Y8D6/nKeq9ZAwO6l2R5iBTyGOjm5DIPMHmqZX7rJGYIl5BfZUjbtGSZbTHD2rqAz
QW53VRMcfzv0IiLzwjZlU9t73ASUfj+IpRXcBktxFxqD9fUSoJAQW4MYdpEao4ES
h0+8MR8A9mIbe75QOL4OyY6P3bD6D0fb4cQxMv7S3+jFtXteQXmaczxVJQvaU8Ln
xP0FxMKBF6XOLG43J1QT33x3wzr2u/BLIvrX94FSIWvWaCizdkE0ZaIh2U7mJVyO
EyXYmCwGFZPOuhXtz6HC7Vec73DdG0oxxRmCDUvsMVUj8CWN/JTeODfaws0lAEiH
UhvnqsyTK+HmT73A1RbtgopauwRl/DRkRBoS6fMhhdUw1axAj617u8wuCKmhUlOD
c/52plx4Pp+bSJQMBP2OZvUV3u2tjK2DPb1lv1rYLcINGTtvlF0BwxCek0npmXXs
Pwegrk8q3t9CK5SqrUkFHF68JyGm3Yn9vefGpxEh1Ew7/q0kZZhiMpNy9Zt9luAv
Qyr8OkuCsBD7e6kV1ek8vmPaPFe5XstWi1HFyZqsB/oXV97z5gsb5GDHhE7EfMdN
nirp4nESs2IeeKns5rgP2jQW8wUrXQcv7PotTV35L86GRxaW3jIYHV8Wm4Pt9GOP
VhcHOtlq/98ynE6yw+TdZdviqIqByv/IM//hWvD/WjuC0oMr6GoLTn+O9dpeucbe
hsbRB8B4A7qZuJQJ2OUsIbpdUQvSQ3IeCTnbJ9iN/lqPYFRnXwHiDNppmkvqOcwn
DUGkhbnUs6GAvibNiXayD5ILUIosvlG1z4ja3KwS07O5QusIcU9xD8G8M1ebm/Cu
HeNSiMV7Q6SMOUCMmgN3pv7742C3l9YZbopgPPLz+US0s4xc81wRydDw7sofP6QX
JqFYhfbWGXp0CU+2Jez/Gt/Ghh9Tq04X5pRS7V4wWsg8mNnTb+8Jbe9zJWsVFBZm
mDcHHsY8IVw/1kqPnoQJVC/9xn4giL5Q81Xox3ISMwEqau4Nig0X+P9qzXbLLpOp
TfOBfeeu+gKQWgRsvX7VBWX0nbdTH0hLIGcl/BGkaBMxlhxpVcPeqK4rlJm4MQza
LuUG1fXgJ4zHVsAkPd4tx4DCiZBmsrj7I5bRmGHqvgDGaid02n9Jdo5JtlkBRoPE
BmYzobepJWcG4o/r/QV7CqYgRX57yp8wdaW/Pav1qrRo+WEKTmeWeL18sUWv+/dx
TPR3rzJ4QGGGl3+ODHUCqkUXnC0MuKpkRdHQ+f9nEiLxd9nFsKLb/HTehFE3hLvk
dF1Vk/qurloaz7ON/J4CgeG4dEQqpbKOasOkOh4dCAitSDAfc6qhPrqiDOEzsgUi
u4D2Kg7S/UGmYWrYB5TVnY+EO3BWE/lTa4/FEYETEGuM6QFWxSpAV9BiiSt0iMDD
yz3kscd6jPY9V1dxXGyHxAk+uifYTQuH337ZcQztXqaAu9qm8L0nzQFbDtxVtBRJ
WsrQpgsJU/3IuX5C89GRnCKC4Y/c/G5NsFy0ehPfOcYkayFIDR0kQUjY/qXLT0u0
ALnA0YSNVMAKHlueunN7qnUmU6K25kuekj/dkdj0ZKMVSOvTu41EhMq7JhpqXDQ0
pBT1ScIet8J0yK9/c5TLUNLyHJ5TjLGn+7YCZVykCxveT2iGEyRClUZF2JUO2Knt
dj6lvNozpmkN6cYmkWJH23JdvGVfuJdxjn9CrQ2K9I0rXVQJa3FqlnwkjT4wfDuZ
6fejWCXb6C8Rpz49SXuRGYzIxnWwuyZSp/srbUd8pX2kfNx4DGStYco+Vc082TRF
OOHammfrtjPEyh4Zdg9uXsHRYdnaObfyCtNClIKO96Qc+HpZ1d2emeuDdX0DkdRT
RUOzfIa0lPjvAMNhHlGrSCxz4i7/7JmkaXttn5lcT/krGqEZybR0z4FzE0SsZnLo
4l1y4FJekjjpwo6mdNLssDzU0v2qwU3piDPD6aVZDzajzZ9T3m5ulZPixA98fyA8
zMu/ZYHZ4kGC+ZtprSjEiaI5teXp5KivtZVcdKVW9NKrTwaSjxpkucEK374pf9s1
FbeTcdO4ETCxW/3ag+RdeOx4QzVceae2Gs4l9mzD9d5opwOkuQsDBMYGb2czi3Qp
PNbE/rk8DTKJXbiyRP80MUVEOxbQ/YIupSVZDhQR5yFwjhSXoAEt9Wt9pDjZuueH
C73QIvvpYdA+UuwgrmKD8tfkLncn9NMpkn069+MppcQQpLyHeP/R2C5JjFjwPHuN
vJfp0MmPLC+9lSinyYtehyEbROrhsgcwhjEuOEVZNC/wwNbKRhONNEkvEm1Bj1In
cWjtpGARuR8zcttgg0QsNIqHdpoyluESpxWvl+Ig5sLoccjMJg3gM6qBQYGgpm10
PV0w4YJ+/NrYtoPReuSGxcy3HoTuuNU6vo2SIbCPFRzLVVg3KmEqG26jJ0ymXPyX
aFm9o8mGhhPg9IV7aWmCrPeXODsrgyXtPic7etVlUR6i3kqCf18LnaUgpQRH1xtd
+2293WrOCcMhW1/LbOvb3tH1WMxiyTLqtG25uPd+xK8SuU1PHHIegUlHhOWldEfc
nkMwGXsLoJQoloUUUGD97xb7rHsD7yawHI2+RQ9SjqRzrSeJYWio7knh7nO+LLB3
07pxGuRR+A+r4CJSshudrDmEQHIt3tQebhwY13mhwy8qSF6TRGcUzbFw9/bZQzjU
7x4+eMqWp39v1tN77ZAUWprpI3eTGrko2Ysf/NSiFfT0QfD5yXgOWvIyf6lScRLQ
r7YfGIBvtOxyOEWp5Sj+/REErQ6rYQF6a+sZOk9DDT+kqe1/W4SxtlH8oqB6upz4
EkMaHqtwh6WY2jJSzoY2MlwTsUlwHDr/1owPWz0S7sgVZsUD0JD7Tk+uNuPkxlvn
bnyfZzijvdcEULOMM/pdaa0ynly92winpc5We0nxFwbsWT1XtAZDOx4QRabtV/02
Y1sjQmlE8aJWhnMNZ/pAaOKOxX0Dy7lvEtmhbzsdTIGiISaJ+OX6ooJehoUgiXO5
G9uyYj97JKkHC8B3rwfurfrLr10aabhxIc6jWqjkdBjMQYc929ALflmVfrpqsDab
KxIhr7bmkPgdcInGDwVgJzvyZwnLGNH7AA5IHzjINSxS0IUHcJS6aThvCeIdzARF
kVtUFTygK6XBuQbiZf2Aqe2SVoIM5XZKXGMHkSXR5mA9LAJG28zPmZ/as4NTK2BY
paZmUor73wKdxwIn82ZXkENXW0SIWWpdbv6JiiTusvjVmrqJ4zraJPIRaQjSgbRu
H5mMkhOmWY8faCYBtrnDKE3TiJXvMAR0ZBpfM+tTmO05yfl8NYbByE3pCnHN7eks
YNR3pincfRvNHoT6ffCdRBuqoDePhloDABDdpF+8v0MVzVhj+Q4/sXiVG7AvZy98
MitpIblcolr0PN7iPc2fH+Cde4269f3qxPCCcYlQMhMrG8u8dzyqVC3D7ZsyNKPe
7CsFnldmI4xmX07S3O6CPLKXhEZaTHcr9bq3N3b9Zf0oJuM1H9pr8+YRBv5Re3na
InPJHZvpqcE/wO1JcFDvf6KI1QrFbBLs0/ezob6WAyFnE2cpcn95Xe0HEbUOtSVP
07jxIlralrlyKiULkm+3PPbYqRs+c5kJqebrfJXms6TxQWV8M82I8L6gLXjUMDXZ
aFFp/Oy3ixivsAjpamHaD1YnSH+oy3NqV5eNagAlCdmJW5SlMyXfrGsoA7JyHudO
hOUwuze9YU6UZKrVVfHH5ZbdLS6tBU6DuWfWBu4qXX+oP6u8Ely+WFOqoZrxMM1M
zNpNnKAbi8v/sOp7PNvKo/Cz35iVMOlayxlkTY22J+KJxBaEP+ORBCXy5Bzg0aph
LMRfhTJhos4ctgxdfuPaO3yRIkTdwBZAeFRHN0ozTJ3gnDt/nTjI2rjByD5LF3en
o2cHJ/hcEhZkgDRrl9GZnD8JxH2jqPEKSONO2CX27tiL2SDrNvp/wKiLu2uoL8mW
DOYC7EdWqAOxMWOKhOFh9qM34FyM41btT/+FTI+MGW4rOJ0yZNuV9xGy/HY9h9Lb
mY57PrIthIXMWVn6ozsyXmQ1dsnI6ON7K3kY7DqHTYvyOZ6oechFoWb741oQ8euD
HTQlKlHzzX5lo1JqhOr2xcfpcAZR5L98YfmUj6hJrR1oatG1qjy1QKLmZaRJwM1T
hSixUQIhLJYY769C6JHQNVPnyeVTw7ZhiW59J72IJVF9dndbG5djYlzzj4HsFwZK
PQmoNbr2wqe7Jt2pR/JmKstvvVzGKv9MmOti3o8XegQcVkz9FYTQbTXuKKpxTGMQ
HojG/Qzvp44nGQAKR/pT5WMOlvIwD+5X8oGkI+rph56M4I1FvEqSvIdhpJvbaC6D
TH9fmHVC2xa2D5gHxkjAVfDJnp2A1IaAP6zZI79CxyFnUvOGnfrC5zdvzZ3Za4LE
jaNAcazoCnOvyz65Zj0DWPbbyAaCU+cUcIyVqpqwkl6825Fz3crMA2m5MNJyOr8J
OENUc+jOIy+CQ7CMuQSAQ5059kUbjH/kKzw1qX1qC43ED2W8w92RjjVCjmTtXtHV
oEvoUVjuxufFxgAWMVybbfj9/8//vGHZGT/zwd5OvzzjCkItNQABfWEYvYT/SLvO
vtYqMwSdSMx3xsUBwbYox2SyjeoD0Ub5y6ruap8XyNZJ0NDnsAPyAe0HSS6gjt9I
TMp8l/aofo1ajARL0pf1+5OHRokN2yKmRcOiQOX/UVA5G8Mhor/Y4aBKpkuQoGb9
+ym88r2potOYw358bnDHyP1XlUEbi8tMilHCmoUMQNTTUrqLoWS/Tr+IsArfFNFN
dH4MqfBwQKCSXVjQbChjPxYDA78b3KPAOPbIbV/L7RSB/qg/uW+WSpyuUHpAItRE
4UEcJNKA/5RECieJ/ZxEX5SqxCThTpYEzYHUtAWM5kThrfgS2WBuOnI6A0Ogc+c8
jhB9akid/QkHilu6x87VvrjUYf1lXB2LRxwYodR3VtQ3r2LxaqnISMPfl3Uy0d3I
ARPGc89TVpUwHkHCBeslB1BxRt6CSwopl0EvtTQEE+xCweGcVLMOSLD5TteBfJp3
X8oXS1i99lVrjABsW9R3q3uzluGx0YWIxOGOsUTWfahno3fbuRIiZvmjjZLI+BFM
xa88tUGPS3AbqcZJmrPIXgSzZneSHbWkHCJwJCrVTvKUIWHxN5FtDT8qvW+ZNpSQ
iuOi7Y9BPX+AEVZua4DZOglbd5NQT7WtNNyC1KNsa0O8T8hn6AYXiVUsfaAWawwA
3PGUoVGD33Az0fRNn9XQ12VHkHPkpobqhKSICFAXCLJiaZbSMvYItVMLRvJIBW1K
2Hdplk0WDBoV0NWNI8C/BMth7HLDSo9Q6NEfzkGv9B2tbSD3uChnkKtOeONgKcPx
3122zAasHeIdi8bLQXX26t/y5dMkaMCMFmePDfNY3JoAD/FA1krDZuW3ZIMxzQYA
QtYpm1gDVCJ74hLlD6Ejm9x0gToQkXrWZ5OBM8Z3dxyrufQKPIIihqpOIFcSznqy
5Tu6hsvZtx6B9LgyVgynkqpBOTVzt5VZi+l7yAPmbfWP38ln2v+kJeGW37KGL8RZ
ajV/vLbJRxass8qZ0GLb2DchM+qA0DcyL8yCnqUyOAoEX58UBaJHKPpJoEUhr8RO
Kk6NP+uJw+hD81t3KI/XFP/YOW+/Wwa2l4yruzPRzRPkv8KZt2XCLs0B4FCNGnKQ
LrkeFHZV/hjzERWy34DfVe0zBIA5xzDYHz8ImQ7IuEPjhLgsEyP/NJ4nbBW9/5+p
AnPWfF8BFpCnugecRaxkHOO8CzPp2yiLN0aaN7CBVnmufGszOxsceCl6JEKLo1ap
5Mw/kW3T2hrn3TNrIbh2/h/qeDmG0VcAlNN1pOULRcryJS/8c8WMR4QVYWYrQlk5
Izuids+x9lzbxvW/P/o/iWFIjuQ96QdCiwY5TQtPoi58/Pefb1vOI+bZx3fO/H01
BbxYXP8rHXiV4xinkQLn5Gd/pmd/b+H4OP8Ql46vWE3mWMPZbYfc13Wh3pASbBg6
1bbT9Yx6/2NAq60EahP5dr4Zf8a2fflzze+qaefXorzmW1H3LtJm5UUVcTxAfgLb
Ib2uCzzoGhYZ0otLonhhN6AAe4BeDJRcuWg93hZ99LufvI+z8oTq4NBjmUK0V+tT
DwuvO4f/6d5gSlWYiiJ2XRtgp/cM3k8O8kMHeCTkF8p3lICzm/dlMjw6Mc1DY11K
qqitu2/yDcC5kWv44qs3Yywjl6CvI9atKytywl4zqNsPPMUicZ+XoDnzZh+63XSR
yJuPX/YrVt7JQgCe1IbrQbCPciDk11IYGXu7QqH2Jdg/ernjD9M6QPJK96f+fpLC
qTCPC7PrpQfVVc7CUFVqyaBMwjAdav7EWoKJ9pnydSbyOpti/S/Vda6TPx7fSnrM
EQnNXCmgBKffbucs1dhZBQHxqiwBsm6NqzPaydwtrBETYd5ZZHIXYNMN2Q3NT9p1
86mN6CgTp9DkJarB3EnZEcgNPQ+w6Ed3lf6SH1HL+hBeEmpzUbXzFmt4Y3RV+3Cq
wNEhoRDRMguMAK8suTZYpFcudg5f7eFSxac9cC/VdEF1QFNEDuSIaGr5ByX+5lRm
7GlQ0qfbbrK2OaQx8BpTWf3eJ87SoTFe0aK7OzS3ULkJ2BdGdkk0hkH1oMhDTdJY
V8hqhxvFtd6lqBQwcdIse7HcjOAEpzdhwPY4i82qbt19irG5J+b7b29BL/XCftVp
0yRcj/w+/41B7hx5mV4D3mQRn6kOCjh8zfzU3alCAwloCxDVf5WjMLDWzXiKJ/dW
QZIx8HJdIjanPwGdBEgRPIR/14gbJE/bS96k+bzu+HJva2UEesjD4Wawm2MV/lL2
R3Nev5avOBCxMr9hZ1LZER7kGlkEBR1dqIbgYNkZarZHOpkqoryM7v/w9a45tT3e
D51s7mwEC34W+YClbO0xw0KHcuTYFxW+ZWagOtsbnWM65iDSMcNrHEcy0ay9Y4Qy
Xb2uve0u/mPG2noJCqny4MQs+9JeHoyQouQB0q2gTcTAY1q7vVddaOK6f9IDJwgk
jsvSsyZx0/J4sO/BlOcOtvysGulewtqSj3CM7mm2zM9z3PYkACMTlHccN1DCULfi
D+4aBhPDxmIKQjbR1fBxdUhctf9JDV3ovkPSm9xi+6QqSTkVi91imMmIXga4LYS5
j7e9spZek8m+PWPCLJ6Niy0tmwibhPC881P9o89YOOX0YJlOdEUY9jaMQaaKPASR
Inny1+ck+fjFZb9oehnZKlCiQcb6/MonV8iVYpaWjvZMtowK1TK6cGb/ymp/AdtW
Z0Wi+46fi1pTLL52P1i1Kw739MK7IkLIPob7H5qgWRiX3KyDFY0H1kOpbBHs6LsZ
t+ESybCJlYBPwpEp9jJGGXVasxWZi4kwzOfRvAZa5a7Ifzts5albtYi+6TY19v5U
4WR00AGBxbLrif1U2/PpFS8+XXcNhIRNbmCTjcbB8dvUhIowOtO98xaNvrFciihs
6vzlS6UzLakpNHTyBW0sxtB9VLm2LOYmTSAcOJ7kL6PxH4zxffjLi5wH+nrFYyHd
2JCKgDsF5QDKdzNW2giyx7dZPk4wc//OSi+EQ7/9eln+8/z4AeEY3UrbMzKlq/1P
TDZTOVZlEQl75pWqzAfINRLmmjGVhnbCghNFf/8xtVvlbfxgjstWk5LKN8K4tXgA
bXktRM9rDDRd5gyAmxpmBRUuwc96ET6qT18ehk9xWw07YsCu424GpMuY41hEar43
t7SzlEalMGfe/DcRG2HaXuVZNGrkzBCQ6NCu89CUIG1Wi4nl1lBLUn/5T3gQTnFL
lCQFvURoKgrsVj0f25EOmVb0sDGMYl5y1SewhwVtObuTK7ptRnd7Te23JKneAXw0
GFTjD/LbfzEBsakX9UdkAkR8Bbdeyfy9EOIMLmILo0sNFoLvvO0lQqZESAGOqL8z
O9EYRIEULXDGgBIZipraFi3fHmiLf8H1lzQtVr2c3x/ZlvdcSXu6PvaRi0UTi4sb
qNgCbXZlOtBRqdkKGykWNroieizTB/OdwyRe+ImrYGPKONc5X7B0cPYTAsVGZfJ8
EiBuO80XsYRsQM8YrCG9pCJ8IfWPBMyMkilZs1U/Vh0ez7maQXG7NQErQiv6SSP+
9FziyKT6Ynd5D3JluAwD7KwkVPNCbthCy9PKvuqn2GD8BpEMerB760QptMdly46Y
s4qGXMgbpV96cNWO2uPJAqX9Z3UfdsmmONzG0/CrXL/u0ChqlnexEwj+ME/zgHBe
cT+kmbmBhxO77hQGSsaRYwVZWFsDGyR23fKZHfBed0Rf9VIYuDsLxClZdH68DDcB
FZ4mLnhmUz1JN2B9xuUk/tNxSAAA1C2T8eWqft1eJ2ul10wV9RElTiyM/MticlST
gPQP18TYikrLsdTv9qABgo9X9D5VDtEBZmqGchPBO9vQX39T191Xl6LpqZUSPE41
S5TRjk/Re/wmsFGR/aoICcz7NRmQVI38DJ+TZIHajjaguZHPTJHUptPz41agRloM
mCgoxckNidoF/onOuse0w1vU9oqqvA1zI/iHhYCvJMFmsBcaanhjps782BFUaK1V
RQuLfBtACj4DG04iz1jsN0p/F/RhqhyZQGJNqAS4mQI0WsU5Rqp13DbguyITxc1P
yTGovGeqwdwLghqOJrWG3pmorVMTC60vpe73PNELjZYSwfbie81OyzKv5GVUNIQF
hKcK0fAbJ9K+0nqrmIwjJ2rtLS4hr7dyVgFEOsRnCFrHR74MTUwUSEyH3tiPeq30
q3sJQ/Mt34UQIEwqQFlPfllZelk+YIG2d9oAWpSAsTu/Ic8gBNfI4eIrrtg9wAXG
69ZqE6fFNqRrw/+/AkHBTc9KWmBCsfnoUmsKDHE0gfbYY/xW3ZVmknQ9KKyZYnno
fIsZs9Z242jv0S2N5RRnP9FTbk7jY7E4JCdc++3ucEp9nYj5wGtQ77usXwGGjlEa
VdV8c/JEsfG4KazxLZ9pouNJe9xzagCIuLUILAxna+M6N//ykiSoSEPNNsDiqhTt
tva4dzBteXDHrQd3hdc8dFF6Na9LgrjTJUtEhg4xQL2ZbbXErfHO71jV0oADfOVf
v9L3SuHub5ztcafBDChGlWaJV2NQnr8TgS6glfo3iuXLIzbiKmuEJ1dHVftT2JkZ
dbKv9SXjTekzAMv9syjRnDYFDE29aLQfC2Ovrp7V9jh/O19lunicNdlFNP3W78VU
UH3fbpfl3ZgWL49YeLf4S9Mmjzfbn7UtbnvSnDUoJQzHtzz8O7MIjkThte7F1wvP
/Ue5CkenkjU+D8WJtqVq2Md2N14n4k2n3JHcfJFH/yZcjaGP1NDPclHJNbAP8/H+
LRCwrOPlIUOSTLAQHj35sBG87DxGyf8t0gw3i+m6y7BmytIhVdveJHrWkt56LUxC
8IHoxbyUrug2ILG1faVm2LgmGERshr4SEtZ94rry68DZhip3gNWaeBnrT2T8NpBj
8LlvI/WSqU5QuIlO5D+U27LGY1VSvkuRLNromMMF8hb2cWJShZXM4tiUA/IPDyco
muqd9MnpUqAKWMFRJoD1St2v5VlIhHsY3M1vNVBZYTB7aCv8Jr01A46QHcWW1Cke
+wNlL51XxtkHdz9kDpN4jdWzcwgYWcihqNiNLe5ocjrBA/Xy6RlU7SdVt01ua4qZ
6yHy7+DVB7/r3sZqi5OI1CnSh7S7irLTcThlon2mnrxBomgUoEa9hN6VCqGkLieM
bsHY5S/B2+janM0RIneEhX36nWt/0lV88lIw8s4F1ku6mF1glr9Q9P5bEiMr1FRb
+LyWpH0Bortutboq3e5iJ6zCU/EoUagzjEiq0U52F5SpvxJiMiVZJqbVHfqiRbfP
zcf+5hs2hg30dWYOUD3gknnd7Vi0+tfI8UQc+OSvxbEac5aCjYiaHMEFd/GqiGd+
AphXDjl5UuYGdDgDfqGwVSTcO7zJkTZY1JQc6ZbyZrBMj42FEIuqrdhJTdgLzHhH
ogYQSqQsCT9RM4X1w9jJG5KsGzZEkXyj6vDDQeCFqfXA5QWlOAGSAIvJ+ASoV3wK
BKAnNa64zUHt6jqjq9SDrsvyF8qNAOdOispf+23tLOmyUXs7wZIDkKEAU5jukewI
snVBI/UzY57yDIFMo96Tn1Ap7m+/VHORfByN/Xwt1pha0+10Sie3xu/XmzRMRGS1
eOnjC6u0BepYhmG9poizDa5Ieufd2q6Vbyh2r921Gbv15x07E6oGGNcKOGPnADbE
7JNbRDlrM5l/FG7h22S7B3GJ6ZaMARFPlzllyh07O4uXbDlomsN7RTG3Fk0iPujN
//dbyinpvco9uaI9lOGqy1BFfs5YgyGM4J2wHJRqhQpO9dQ5tE5ImYRLYcV79dl7
xeZ84pGoT9qiWOTHqgHPA6P6/QADLkVl9NI1MLg0D7EI1v9SXclSQf2EyxwBQjad
B0yqlaFSY13Wy8wtJzpY0Q6DJZLQvpmHINWxuKDfxo9KRVeHkLPOR3TTkpiM8OxG
piW/Hcf7NQtzjQg9fOE/AAqEsSwkazmeRCvNVUw4rlB6e4T3kimbNjSNlXMXguJv
v5pFqdw3KwSwDgLwHyZRa048kXb8MpL6exCPQU1HxmZrjX6eRq3Gapf2OT96+MvF
utgsHOhMk2uIc1wnFg0Z+K1w4xEQz//PnxplulNibAoOFK1M9FqC4Djokyfvqod8
zLPJqF7X0I5vK9+S9qAlPXoMRhMWnFlghrSPM1weWDXL2/HUYRFm1cmFS883mkPw
Ug1abL+RWIQgAFqjRdteuUTPY9pTlmrAeFvKIkSYH6CexB6iXqj2AEh75fmHSp0X
7blICXq59vDFx2gwmbXWe04IE2HmP2FytFPfaZRAZ3fwumYkxDj3ldFbZBAF44yf
4xNg+ImNDa0oXyzz17OhfBUQHpiLZ6tSumh7Xm1NHcEqdhG+1FxsdciNErYj1LZE
kSGvrCRs/7rMOxTvGQAab//5bibH7Y2QSeEe/N8w6bJYjsw4DlTo+HyB8EEQ5162
M3l3lUxG/i4ta4tWkE8Vkdg8P+hlCw02mhbg6a1SFcvFab4x9QoiFeyHbDCZ4bJn
VePYWiCwPbkb0pjrBvMSbZZPKsDszHNi5z/cce2GlCUxsWnvX9WIfyGf7EsZCc0c
rpnVuqFos45pVjppihDhJvvD9Y13vxF7SS6bnjQJB22jFevukDlECbQgodNeexYl
BSMZOcva4pEyuBCnBLuns9vMc04PJx6J1YOxFDhD4OjLjDUC9Y98kkTKykkvsoK0
Y35G8fbT8fCjkttVMOtzBrV8rjroZo4DGi3yWCmKc4cHQtnw93S0H5BfdGERd03G
5ZdwBSreyrsm6l3p08TCAdYgqkdwCL0bQ7DUGjxYMmZMO6FhwfyePQ8vUgtJWAv/
cS/Heu4ZkgEZrhH6AGHV4yzRGCLS4GICImVkmPNwDs/rwM7jCiNjE1tdlRqXcSR1
P0tKaG21PyRSdE1cHF2kYrOwfm3skHuupps+mWR7f1fA946njq5wLVAKSzGmNmgx
wqU2AwhBw3M+5gNwPAWjYT6p140htTs5BUeFM+8KVOHARKMAMzTht2Cw5UxD9c+f
Zi8WtxjFzoe1GbNwN+3wqjaFPTXf53hsw8+ZeZPVMfJqNIl1lW163T1GmzORuEd9
jQuk+/jvdW1m4viM0VsIqr8Z4jQh1ZJeEdIa0XXOZUaa7ZR7hGfRg956n9SlDTDP
RP5fhOZwCwZh16C8L05ypOeDvMgAMfeWuLkoAMEJlcWvT0qDe7+iX08M0XrRp5zi
25c7G/Jh9XKOaaqbkAN3sPKX46JfFB5yNksnc7MgnblhQcnIEx1Arp1RkzteZwTc
hTHaP5sacs1sizkG60mO8CdVJd9F1y6PPw70p4VhFJ1GlcL/1xnbFl4lGjuvXXyO
QI0g7TbCcYV4ehqDtFHA2B/gbQcvFUQcj/iDS4yLO5PWRhpgtM2yGuO4SE12oIRY
UhFNYPt6uGq3vgYV6CSjlI6L8s7W3zMnhVGK+lbxeTgsfJ6XyCDIIU1Eol5Cr82z
7Y+UI0ekBssHqtyL1A6Zb5dFKlnAk2tYQ10NBayOOIEctlwTZ6y9aTscim/ambXe
3oAQketmUqs3WLvWTMlhbDsQDCZnCaT1rCTqv0tipK0D702HhJwGl3JnQeSTEkGL
VuEDD7WMVIyWgSBWihiE4my7Gsh75cyoi4DAsjaEOim1LU8suHzs2bSKe5r8D9RH
II9OzCMjKN5VoWzufZDcJ1BFhkyJ/of2Kpbgup9VUdpDewj9N2i+aEA3s61IHI4F
qpZXyEEy9cYuRuOLFhNgZSge9WPYrsAZU5EUYzE8NjnSNJg3XIFT3Uzburw8fH0M
2mBXqJ6jprkzR/mIOwfN4bkYTrWVk+TvrDZ4vOxkaKRBCBXUXc3p8oRJ1kqGQ9bj
Ryi4iDfyRLorYLycN620M6lPjXORYUg5N6fE+EcK+IRSFnNuJgbAnbI93Pevs3I7
g5mcJRKKRlRP1DvFKzHSJN083rtn0uCqlUwcuij0s+3q2uJYTgJQor+V+yK8NHJ+
x+QzJzhG9E8i1f0Ne2+eiESKdfTCtzCkhVXoH0HiuEAtC2gBC2tuaJXzqpGlBuJn
NXLESyNW0P9wTD+1L2qcjpPyKf3dwstGUaUBw+8Nacrbl1r44NuHLlB+6U3ANDNz
RnKS6ep1f1Qk08AicG6YLA02ML+M4i3ilhlyu82TPcqRG54fzIx2zjw+VQGFzTD5
qCwJua8PUKuCtTjtaKO3RmJEQyz8TGWs5jY75qtipgCgekUrgGFD1LvZvTgYjr+i
+WaTpEpgQump3XXt8HcgUerIoigyNRcj0RP0poHoCGtjURjv7vTWKBc6vSKjUbw4
9ql+BhtKZclOQcxsCnAuORSEZ4lumIUv4TWPeE6FgBIj1e0qmTULx+X87ilvFzCR
Ty8hGTMMv3M++9xkWBzYssIPLi3FNGJj0pFpus8bXx6MIWJPwI4VlvS36HBByPZR
Gmbgec1lzfO4EqrsNpoae311GYnvx8xUydJvHdrIJ4LhnXFG8aJ5RypuNxeXEDjX
pHAJbJkhRzJQ95zCJUCSVvzc+Z9B1H6qWU97h9aAPH9motQwSSLbUEGfGvsQT6vC
GgUAgtXO1Rn7T/xRcsumSx14oRriDboqShCALd9ZnwsrKsk3/+vnuCEnIq2+2jLE
4DEiN6W4ecJqRN5kuMM36UpXpDvOzs77JCkMJrXGxbn4OHCU0D7gO6fd4wAZjS/K
R0/Tl7YrSa2Koaz8XiRPnKe0ChYR3JHnYEAFDm5QLncCWjHUL/lPdFtWWv/hRJJC
2HxoblUedmYhxqaVJzDuSrLRcmV9WlYJcb1cvV687291TIjSsjql8efevy8Uya2x
ytcyaMCHti3sPwTyIBhCIBFisQisJbvyNAF+Fe7Glf1LenBvzBOIn1uSNrzbT3hZ
HZp3ICkR/83o8tqHRlEXHMTL5u4+otfseGZjJE5irPEgA6Lbxpwd5h7089rrzjXL
zPeky2k/F4g5KRgdK6duCEYRKwgatdJdHPhAuO/ASTzMslC8yUm0wp75Owxo4KFW
ec/5OEHmXc96Yocafqf2rxEzc+lso3nMdthlnYKskLzrb5a8frd8duKEUDq5mbDO
ofHdI2JunffFDWT/djSjXAPyS6whhO8LERDuPHPXUf1Odx+iT7zD4VkyoQGt6/mu
mX8zO3q4kcVAKP9FfJADUumJn324osnT2/icY/XqKC+eBiDdrTdYddSkFkH9GbcD
HJCI5QLTDdvYsZNQ4EQc2Als714GKNDHSvULzPXD3sAEJQqWpXGtKmIKHEmTjK4H
A8hxcjlFk9kBee+NNfHaPGrtNrg9pNig83/iaDOvKg2ncMQZL85IA+USE3747nPi
8/RcdMbxHZkajiXTZx76LKpahyQtgxxEU9Ie+xf7faLRcXBPPLtpuoGHrGzMXLEJ
mLtCGaJqA73033AAHRdNbCP+UjS0WEitJDeMLWqv4aZdr7z4vGmAYuX+abzZzmIX
hKIXrjAbciaV21eQeL8FzOPtirvvvc6mgspfS4DHLjQi9U8zGrhxLINKrVDJcN/c
q6q5v5rbSmuXXns5ollud6iI7iZ04y+dAwkhSKqd/GRpav7HjVOtRUghwNjji0H+
5lteBrl/e/54INre2VLpMcLFEU4xCD36bh454cRHBTG4k3dUYurs9Fs4FQ07vT25
NbzJ1GFlhAGoOCRkmmBgIrC5umuTz+HwvvdsmwTXIhEvHTevhpuEGMZAtsNGQKtX
XPeFQjU7i9fgSGn4JG0e5trdDhdyXf7FwxofxCdhFyLdFuLEqTJlJaA0OIfzdNLm
tIvUJ13Bvmm0HsQIJXlhmPjiRbRNOrnbIbQMcAxYEi8OZLRQakNdOfJaQALKdU2M
/UGuyTjuK2lE2BCuVZ9Hd+ZbnGJu8lQXTwpHcA9UO2hR+jnY4TWIbrZ89wtcMjfU
+f4Z8xKDUYNCinuZ3SmOEilLfvEtW/ioZW6V3yM25Y5KhVVH4dbaCNP8Oisul7Gp
BWViJ0uzXzu7tQsG5xheBrtXCuXkUC2h9wwkgqFFAvl3Yr0oWu5tE7XYUG1tmkHr
xEXUCbyEp8KYDp1q+5akih48p1L5B+1gHr/HY0cm1uDKDNu8a0UIKkvfQSh7aLz1
o8DMbKGi4f24bbYVwGqN5quq22rxJpUgdf4xncv0WacLHFVtOraZzVwyKZNOK3Ig
N40ldsU9Xb0lr8Sse2I3UJOrR5qyCobKYrv1BLzGa6AQfnF6Xgd4IEqyEOfJQLl5
Y3Wci8m1msVIUALehgDTyFQm+6Fki7VxNongMfMcfhCeB9rYSSPlIw2TSmOaHlW0
0yxix0BSwbzI7XtI0mtIbmybhybGkLwd5VRPtb43+QL3oTiA7Gesx4YNUZR7JaD7
FVFdY72PrRgxjD1kN/SnltxUVEacVy7m2eCbmhK+E1Ign49/wA+FuWyU3nlGTiR5
Ba27t6PWiph2BHYIWbB9d1Cq4jrFtjhsEwSqEFX9lonyCEzJV4W65DDjiN0RwmSr
4XS6tqxIb4lYTGUHFkfqoL7sb6zg2CwkzWrrfn3Q0c6UxwzsIdty0QnK0FmSB2tk
GitlHm4Y9M5SUu/mIs6wv+lYb3SXMmjFmAjFUd98XZEwC6VtziP7IQYdH5PPuOr2
O4xcTzZUyECwNAbbghIS0M5H1Gl8ge1skl/fnGMxIDNF2Vqk8au6F/9jCB4NizoX
ElbCvINO7+J1URY0ifYK32ZRqdQ5oepkx0+CdKFLU4O9TweM8MVyYOrii7ld6yFA
+nQ0ngUt+wQxoBhwnBon0MUq5J91P3/cthhJea9nTRwhN3//Z1fe7vJFlSYISril
N4mf8++of/znSlp5tOhDN9GCSHTzENDm9RYFLPNoFtMR0qeSfgszKuHJx2YtgGja
Q+orxTyH0NNXwX2jc1QKANR0jJAMoKa8zAW79E42h1uvL5jK+IakTi7phQUI8PAj
cJp6w2NAOQnRYDHZ1lU5z8XBW3G5eLlQ4sQ0VJ7/VkVuF/EPS3Cm/OcTnHEjreSC
8h/JaY+tQiIFpO9M22t9+9qT9RfXJLoJWB9SNiL9wIG3CgNK2UnZzmXjwa1G1fPB
kubd6MRzSwfsk5Y3dzG/Bi8rp37kKmfHQD87NCs4dBSoKRFOO796W8EL6ZS29Y3H
4B25N45YVEElOTH0D7gRa62QNE+2y5fCJIsz3z4sG9wg7/nHQGaNEMdQ06EiE5L8
itGp6WIooKGJo6jYK2M5DG9YA1hHXVbEaJdao5lyL/NQdmlYjYZQczMijIKQoSag
q8CWHRKWo1Co52icT24G+CCWIgwrHlNo3QquGrxb6rima22Dkduz3PI0Ba/VuS+D
TbXdbLVTl7sofsVfk1Uz0y4uiUqos2IHnPtcW8Ne6Pl0NTUhuFSvOX5KGNHQz3L7
3mGN+FotsS1m0/TePW3hv8RnWyxzKqqCr7nx8n/FvIJHc8dbJLyRiGJVTjHZ+8Au
r9t431Gfor/4Y7UlHcpTwH4m8nJa6c9e0Oik1PSDAgSSDm7vzaPRGJKbiKKGRSrs
nX4WzyQfnkYUKQjOcGqA5z0eByBdC2Y3Q1IuWo9jLMc6+F6+65Z4FCn9V37XojpS
jZS+hUScXkOv/1XqtyYRwoW4IP3O1bnygfdtuAp5jKTq7Be5EjJa+Nl3gmJ7ATxp
1AHm1rfoRloGbXgKwtGCWknfhGUiQfHsIIdGShUFqV04Vs2s9K3QZ44VZFO05iXF
pKrTjEtP/k1NrKim+bnRbmZelcU3G3mm2x5EqZqIt3rDoISRN+urHbKxHYLjL4AE
rEoGjcvk53U4UGefdwuMjqI2Kho73OuteEl/cpnwxb/vX/7Nz5eRuYv6gpTmFcA2
lJa6WhDlb2ML2yHl7+ISU1icuIfNUXWIZIVEM1FpyxsFp9wz/DPXZm27oNznhZen
9Ns/6CBAn/Dgomb2n2njAEF62DQ7xvOSWYNkFsAgCdqoKqq03JSscmXsQ1rHj7Oj
WY+3Pj3Te8fzj3HBVFD6WYNm+sjuzOpJv6pElRrUNeMyuklAzbLHB4l0Fbp3Z9Z7
7jjkKud1oFu9psNDvV7um+12h1tKoHRfboMWnkhmcT0ZD4m75YRnMt6Pd72AX/2A
mppigC7LqyYdq5T/kc9GSZ56xn1Cd9hcS7urhfqFvK1Iaispi4pVmumYbuDtZSN6
koNT7vsNrJ1c+GwCTGvmsB0XTa0LINT0GdBHRhVNCwoQPLNJMLWIapS0tIEpYjV0
D1XLfP5ISSR6OB6V8PJRNBiak0O6qpbryNyrdIh8+qZ0Wc5fnquPVA8ucJQlzP9q
98qNRviEIguTIcYNXgikMrdZsKUvSb4/20LKkNzlSWDrm457jXTPgRAk2uNJ53u9
q+vE2Ez/L1Gea7RbN0+vwYDGQFUBnvB7SiRC1UoLYAzkSk9iJ4FAoUXoyDamMcDc
+uBFy0kc9cZ2o0QFosgBUahwwtsEw3DC296DD1jE+oL1DcurpwraJibiE5c/VoWs
29UKDIP55AevcU4S6UgUTVUYqGXCymHqU0Ojk4zsphA+cWZVt+5AZ7NA85yqp74Q
LTgoKNXOrP57bqL01OjAmxdvtVXj6f1gCXNT16xMSFAUuAOasrXu0oCdgqFsIsH/
fI4r+skA+vVJskxz5DbQN1M75DXKscsXCSbEozyZHy05O6/5ha9HE/wJq5eUDtHG
/eob9kr5Gtq0KuTcjxoXBROrg2FLVn2WXKPZGIVgotUYrUT+cDDTNEXIVwrWkaR2
cGou56E0+fZkFNoeoyr13/WDGRB8t6+VlSfxET6sr5tOy//oO/1ZQFlhI3C+LtvR
gtvYoRxGSQQxsyNqfYn2dz5r/XJKbCAaFsYotBw5JGCgRKXeenxFR08gZsEwLVzv
I6u/TYi9t2rvH0Rv+zYZTvCH6i1wlg/SUaJZekFM76lHQBqsrMBGJAWqKYeIbjBT
CgbDvJUOP7TmA3w6+QZ0YHC8ABYKPzLd7asNVzUC8nHXKk1PQskm3FECyTjZMpeD
1O3rycU3aup1k8/ASoKHnSX/7ca12DbE0oA8BPyA6YNKHB9RiRC+3vj9lCo/Xoqn
rwdVNnTSmc92EIptwb1mHVN/+8hsl7FgBL/0/byZ1g/jI5nYdG1mlSvKUFu3k4uC
wTY2Af++HxlRjVM8UQDrM3uxgh3xxlXTfmaLyF2114W7qrCSN0Jt5fhpISZHPK5F
AhgjscVwHrXMB7rfuCcBjL23nIdfyyp7J2huFm9ji2PWaNo3Q4OYvCncA08qFYFa
SwFt4HsChM9ujQvWKqrmdxKB36QJEmebta3OsnkxPzirAUeI25yv07yNzr3bfbTa
Q2KjHFzrTf+AQ8OxqDtlnwLcqO8TpvuY5Iuaa42H9pFXOUcHfTAfsh/deNd/WdVA
Jm4uDwxm8BjHt8lTWhhJ6fmuQ1cCmZmXQw2kuoAHsbBDzwTz29qH2/g260QeOOuT
kxFCZcw9Pb41JTVKZCNzaJpq5zKciHjf1qGK+KOQMSihqZglsNWAxfPgij9vyni2
qNRok+Ep+3PszizeLIPE7BIcwDQxhL8F6ptpSFMUBV51fScoph3IFIbjs/AUo4Dh
gXq3GDQruNZNWvCYQiPmBsMx2PgtTOPs+Jyu3ESjsTk1yXjIs0zG5O9LePDnJ/ME
QpJg/AJr1KIFYybDDNigJE8Az2NlKnN7BV9Zo2pvTOu2Wb2AEUlassqshKEyP6ro
Kj2ocwMZUudjoEfLLxGNzTwJdkf8PPv7FUafk0l3G1zNgt5mxnumJvx98j1bZSRA
6CTFBIaBFG8nRUvPRxECrzb/SpCL6LmOvZwpWl880oV7zsZ9TSpPwG/6Ce4yfawL
Fa4IDPnHI7gXzFGNJqKjYW9m5OyguBqy/ZGzNBY0jcZERLJDglGgcp3H4Xz53mns
y/NpZX5lwPALbYYjS4aLpFLpAaMMQ12n3BNhKT1lfBjO7f0S8TzYhIBllo1un5jE
qseCrH9Y0eG82Csz8r7pZDgns568nzrwM21yZqUPuG9EMz648mw24xGyAn8S9zV7
OC9tbQ4uz8iOFQ407nfhjm5gbTI1DGy+6l/BGIl0kRZnp+vRIq2CXyZ5Vtuu5M97
s8SrMZr7NSuTgsuZY8/SO7UUTsrPGKTqHtF57II6D8xfySnLpF6hpE8fDhrI0vb7
S+HzZK2zzyJWBXOE7GAw+TcbTyWF/bQLKuU0l9B28JV5TNNz08whi9KDeQsY2SPI
TlU3DoP3nDQpLEqd2ODcgPpsXem0WssaQUrEtR3vPTDUZ55yJQ8TJX2vb54tk3vY
kbMK+S335uQn7HVtniPIAoiVobecMnAfeZ1qCIT0me0BwCDlKMaXUTL2GAAZyAIM
DInxsBBLU1ITazCI+jQXBlnxQgWXyzYQOFPbWaVBgo6BRlu9CMYCP6BTRav0ugAl
qLGR1g5Po9ATdX0fPBzyNULSl7itgjwQuKyKw8iDwXwM8W6EpDZbhrTmp9Erdqws
D7lg1pfaMPQUWs8JUPgVpUn3bkHvNKI5tCG+c13PF63MuAAPa/Dhl4D6v/ea6DTv
prOTAopF3ggwjoyNIofLPBQjFP5JVrtoP31m0be7JPk7irST/qAX+gLAcowBricJ
2xy+fcMHLquwLzzBCM8svjYWyf24xxq5LjAQu338pW1mlLcuxu+i65w5zwSsNN2B
vsFzJOnyk0wvMgxmlpJ2eiw+iomXJ+3MNV2g0mzlIPvSc4il/ojTHJ93zOcumNfb
dH7HGQ4qs15djADedR6xT6YACfZ5TBcYnKWVNySGj57G2mYRWUKKOh+KKDYARpzv
W/OJ06ygFRN8VOKNzOvyuDGEbSJ3muKcej0wdxVv4jQ4GgimgO7UNkqm/Lm03xwi
8SOZj3yt0+VTALtt2z8BEbCpb60wPZ6cbdWdhLZ2aIRVKdd0CA8quQpCySDOE0KD
R17pWtdWlcl5vxm3Cg6W/bt6NtmW8XlZVDyP4RYknlKqEEM17qs4rNBzskXZiZwx
K5VMC8TPdWaZiutVJfRqhTwBwEdb3YwZnuWW4nIsHNFmvFaJvZuBikvDSR01WSFo
2SWmTYfHRDhyKNaCo5pBpg5dLUeiVi6Dq7ReaYxGf68Jd4a6NzJtyJinMTdOgE+H
ZXiyAvaMHgtvgT3xovaxtiynHpvaFwFf/4j2pFYIBjQJfJi6lUExAMl0FIicaTaa
2+1K7cYfGfINjtVbzEvdUFJyo9UPZ/YvOd3gyIj9X4Md0K7pNYATU7DFVFzHkmPc
WtPNcVowLl/xtb+Q5iIkPBgvv3ZFwGRGOa+iNuzYshV2FEiBHcmnTfTbJJXIfR3X
3YlPgnXQPLDkvljKCtDSxrk4by+tW4AegqO9mNQpUq6pEhLPwcSy3EO81tIjahzG
MrFRibqx3G6ykGc+gbfq7HWV37LxbJ87Ry4srwLxdnAt2cA3tJ17dCod25F53ms8
1SxRaX8jpCN7XjlWZ9SNbozM5lJMOnexxKo2lxGsEXIjEbVm6R8Xyl2jkrLnwcZS
dIjVfKTSSUeQ+htI7QVmwmiCQqvLPH49wPwMjiXlIPTH9ix6IanYJlas/4OJiLSq
BwfQptHENwA1EAyOnMglqz8G5KvZZSZ0Yf/bUKGMElxZA6ODxQqGCYa60snjAKda
CzWTaSbJPoxOXi4bUYjlLcr7HLlUEGdSzQ5cITIeNaViJiN1oPhxgi3/4RnfEIaa
1S98Ayi87msUjXH+xCSlYh7hEBhSeiZgN7GBLaSSxMMb+88LxHK0ty+imt2f3Q6Y
S2wOd+O+uvF+pbyX5ekQPq6G6I1xjNOS4hjF0sSJlMH4ycGPYhbZhS5LxGvyIQEa
eH7raAOMVyrH3wdxJbU0umh0wnODYTXG73QgQXPn5ZAQgsvW3pfCnsHConO4GUU7
mIV1T/PDSwyI+aLNhWkMWs0bG5FCTV9RqMEmK2iYWnpybCO9hzIk0nmqxcHyyORm
004idesS/yRhhqwNZyFfKRPvJEtJSnI8mfqNJ4jS1mG7Q75WQCZ21VInEisSCRky
KzmXhYW4l0WbS8ClF2c0iPAiEeUSdUl3kuKpecCGqBFjFUyTYn5HKYmUDECwlWDP
vPybdhpme30poLCQKjAVpUztlg0ZN5bed/WZJGik3//jeFphh8IoXhw94J13iLar
zNWbjQsZ7AJkBplQYjj0xe7aGGx0jB9g3WIrjAV+gIsfZ5gatwDm4bwSEDVmLvjN
RM3hI6pRYcoyjEPilD1HqCrFJWTS/evC/kIGqJh0s/qnWxSu4YvgMRYaIQTEK3eU
7/3UfvxBj+cFZDJ46jvddJoK5mU4gLIfYGviRgC3nrShuArHEZkXQDY+T1VBgQbr
rfCCKNY2Qe8XzXkfxwSYke/cjfVZJWCL5QO0ufwE9aL+6z8ND68xx2UMLOsZyPX/
/3DGonjaFGp5vMYiegaOhF6U3is80Duqs0SWY6mAAQd4nCI0/510guvyz4UbecRc
xVFIxwLPUM66ClPHcJH4lbFFBVxz6le6mbEKdpnFvysRKaCJ/bwSSWY1ZqQRTG65
lNx9FrQZAQShNVUZ/A/vwJX4RWl+VZf0F5rY1MdKbRRJDe7zB89ujeem8ByRAMIn
KQYcT2/k9FFY8FdluXdQJgTfiSLQXuR1TFxO+7tfeGPLAaRKgoJiDwqLPhinRj9Y
/WTbseveUyegF+0OFhln5inA+M2idkPx2Nvl+L0yQlYppJDP29Z5B5CCq92yAJvm
oF5v06TFdc+zNDufzhZb4AtxzPxCkE6068s4jrwoifwFI7CC9FHUFgEEtzukI7yy
iBEiirI5DQIdhjttQSGyES7tDCvVo4ZnTb12Z7qjRjdkPLXxgHEkaRu021BxLBbW
GIwZq2J5Axxs10Vu0jMUbmeoK57sEwCchxX7zE6N9aoLLDz0EUl7uS7eQdRZblHb
1kJgn4Do4gUpwkKO3AU3VJ5VCKjS8yHqyVLmOpuKc5RguV64+DX/8Ksb9AqeQN7H
wn00n/020hJkq67NPSf3yVSKBBUvkBnVwVJn+XVIyfNzCud7AXjMcF0OfIlQ9UcV
ylgYeo4Nuz6OtgjHUE2LOKPMK/KfPHYmdM8e74RcYXXHu1Cor/OZW1uV2zFz/LNo
9G7P/ykMHLUF69UeU27s6vInmdrkHleL3qDS1lDIALCwsiH9/DFW9r87+ZLL7V5j
poWWzHDtzXqTGC1hJCBkkUVP0Tre7i8LlN5sFH98G/aEApM5sRONdWvMUpUznGju
V2wOkMJaAcxBmS12pmJ0uyTrMvWau5QADMxcW94g5nvVOj+GMUn/oxjP9IEgwXxb
diRtCGlyO1Dg9mYjyZ79KhotQlIHSI/vqlyGGAkQesoe0e3Ck6AT7Ornhdxi01Lx
i56ySSl4wtMpRB+RxQdzvzwsmR79KOdiHUQTt2QNuwaun04vdiR6M1yfb7hdSnLV
fxZ963c8FvgQXju3aN6k3kYtgnf9TnRuV0C1cqyThlj25qIGCRM236pDl2/QLXmU
0R2qfJUzEElZA3o5pJnPEpc/zY81SUkzqWnjPdSj1cu2pvnkaYrI0PQBRfOmgUkD
yeZWdqiWsdMX2DCjxBYNZ8aY53QPOjw/wNJYL/kT2QxOxJbxTzFqMieM5K/l5c16
xs92ocxz+hXMT2BdxRHbcm0A1HwT1xIS/EcIA9x/f2StIMZSkPiYQnMU8wWFY1FM
AvjX8B/tEM4yr7Dkv6dPcrCm/A4ln1PwY9sC+yUwbU/X8ECpjh/PaEJfiUp7Yxdc
2PZhkaBzIL9buu8Lv/bJOW/+EkBy97d0z3z0vjBJwpV4peB87QmtQUNV6VZ2vGzW
maZYmDiHAPvuItNxGdt3H2NglJISE6QSc/fykM70NTb/7LdTqMNK64fTR9RTPM1V
Ui0evrmUFdiK1cV02frXTaVyY1JtKhB1Z3XwcJyPCaDkge/wAOWtXq50fi+GRr5Q
lvd/p1W6qXd08o36ocoU80hSWcrobeQv2vlJTDPcHk1XgIi3b2vXwSPXbkxo69Gm
RT+QJkeDzK2LiZ3Ch9Us/5niCpAenOEq07+T90cRv1zT5TeQIjbkLpj7psfK1xBc
PP7NhQwYmIOoHV6MllxNwbbs67W2AeWUSURjo/kYHqsV/YP4c60Tmf3EQM8wRi0D
EWMs64yFFOuDX7djvmVkt0AtTwzs6c2Z/6nYvVhnrHVOBdYn8NIEr5XddheRCR/d
lmV6Id4t6oW5w7dvBnq4dOygIgy+JfoUOzfmXzXDe75rY5AC90IpYMBFZ6fKzYvH
aIMnxggeEn+Q01fMFWtMDRvATC0Ep/xugw7+QlgjGEp/rPywMZCxA+Vaa6jGFz25
+T+NUNVUEUaI0ENLbxtkDXhXs3EZcixHAwGEWimIAvPCUnsTYdJxmSeE31/nT4a7
5PK7P45uxwVsz0qwnhFbE6MT/Vzlo8p52vu3raYgUoKC5wk5CcybbqAwGAr8JOqq
eFFXqpBJ4wem0HM+D4FetOGzSzl+m6rtFYCS/65QdCrBOXJUbmlzzkflV/rQeHXQ
CdVe7jCjz9AnrwedYbItgJcLhGPvLgdLeEAr233BzEqamjH5zgFjSt993PLLGYH7
ytLpLswvqM3/GzG1/lTPzcWZD7qF43s8OogVPboXWe6ImEGDQyq9sFsC+FttB4qr
KydeoCtcNrIh4SGO2t2XFBbGAXeEBaYWKnsiLMZpdOJHenltlKCGxHIzAtOc1X68
x5illgMYEfRet2v9xoWVs76YZ4l0lBxRT+pVYY4xngEEX8cQghwrvs7fqJkAj1i9
3bliTL3px04/VSgq7Ny4+OaYyax8mdeD0tZlZqsoz8kWDRooZtDoq9nvT0qVtPkd
2ebLrJlg1hGA+9NnqvwIQxAdFjTw+vQKxn3jfls+tFZ3VYIAO/rfsSGvWD3O8Y7/
ZnnfsRSTu2ZXVowtMg8O2DhYQKWGMm9XCM0Ri2YDgy9SsFpbMDWsQoRQdzyil0Bf
ccATRDR0hg9dj1I9DmE5apo7ewY4F/064Kntb3gTun9TzRYxMMfPlw/1ltFGrYWg
oeBk7q05Y2fdGwNpaNDS7CkNweXHwWDlCJj2uJXoWAS3K9h8Bwd8iLw3zUw1KR7X
dQ+jFUTSzOfpY5AuRnzk5p5yvBtn4NdENMStOwsvwKxI0V3cbHyugBkUa8WWfmqj
w5OWrVxh0bzkXxMfx4L3ABzHi8BLncq77OuVBdWnHNXc35JO+vJYr1+G1X0Y/CYX
8J2ehUaa8weIqjN1E71NnS2K/be1ESHhxndTAmcEQQ6z8Mkn3YChtT5JgA5uxceD
SCIY6tqZjDRIiYEv61KUZ8oEACN3ZLwbp4b+UBqhmZh5PAn4xDa4WYlYLdyCPqx6
Sw3WhKaQdXKXN80A1VY+g2kscoiU6yr40zIrsgEEyMYlJsqErOBUUH13YfVMtxAX
DkWyJ13OjUXfmb0622JgHJzEBssF7kolZYix1v/6u90QSEqasaXuNZ5aZphDs+lV
kLKSJn/YLjiRzeB+QMo9K6UwjgsPhSgdvB1S3hxmGuPpKjfFAH8ScfKus9+mci+/
nzaR4Ab51D2IvnSBASX+Ipb07xtKajZMthfCIdM10mfQNhiKjv0hywzWj8ruE4Ff
iTMWpaMzvxqGdSq03tVH53sxSzs9DriMGmmXxB15tAlKCwONBiYIccKRJUyLlarh
OnxhyStT1ipAwHHEI/AvZ958k/+6xtFkeYy3tLFjkZifEV58SDSl8zRWt3cuuSyM
Dq6m/CmM8LD7jA2Oxhj/im0emo9YmmbZ4cLIVC4fN1LDSdaS5cd9eyaxN8r9c9Co
nHRZiyz5AUfygIQa0G4GLeCUNJf8GOdMMO1Fpv8STS4sptCsMEaJvU7Zj80uJ2C9
CCJxdVWqBD5HLirWX6iHEskc5UtPO7q/tNrqIXD9RqQwySsKl1sYhYt59pO8dRqS
+SRUIhcaDv3aS1FRG0QQAX45MyDhlxt+L5MXGNgGqQiOZuDvUbz6dbfLdxUBbPQ3
b5HKeW8xfhqcmfcPj6CsIjC2GEx/YpF4HIe3JCjArFn2xrUBeLvNicdrK1aCp7Yp
bQ2rCG0MWicJOR+MCGPVUA5Uat0uKGEn1HWgqzBxsnr9rGIkqZzyxMpkXk13OxX0
xYJ0NXJQ7hPBoDwcBg/QZqsdCfRR0/f6nUCZcmRfD4/4Q8v3vqXJKG3DjGzchRJQ
ZOs6UlhlQKbzZ2E2p7ISjQJK6IDEgzkR/lG6/jXJDWO7MYcfANbS6DPXi4BoCEkv
gK7Eg92oU9ySPFtEUbWh874UUF9k/r6GiG/q7bO4atfNhXxpAQHY4d/xsgHicljZ
epbFMKkhMZGFn0IEyGDM0rGD5fgPc7e+R121he7JScTVQrbrGCKgKDRF7KXqv5nb
honWbsfx/Mzb8KtNIhZIUHzJYV6pBsHRZdUTv/xO0aLPYyxPeylVQU2FuljMe1K2
KShrSChpx8uzXE5byV4mbV6oBlxGRALzX9RoPBnAlV+j6nuSAjstyGYs7agSl0VA
HUxo2aRNg1+6fi/QAk6cWeq2mNwtObYaHrUjdQmc56FvajZ0NYqwHd6iJOzoR1OH
IjsewDNCFIhBv7irKsUZBSfcRs8ofhNkpnN1x/aEBHe4itTUuO8sBKmO4yskq251
MuFkceI6qMRtvGYeW7617VpfexU+1IoWEiYHgqB7eFVlGcMPNBSAnBjAx2hWKDyZ
IinQGL4W4xMRe0tzEBj+3XlJ+c714mZTrEJwvbbwOj8mLNPrdGuezbj0LjiEVgEG
nnFV16htJ8Hch4nwEWmMWatU914DJs4OpCkPTkUvYtk+YZp87MhCac7cFVQ8A29+
KGE6VN0HUz83GzsJ1hNvqdP5Kisy9pxALWMkBHkzgbIA64vi8xoBsdTTTdQoIpAz
bClWOcgcJQPoYOavsTzlXsiyAf0r+UpiAmVs7BPuT6OWsAWRYxL8IeO4k/+HvnRY
0rJTJPFsZCQAFOSNo4WUgYfq+zvnolo3u7U4eM53+sMt8uZUkmeOojBkaUWRyK5M
CiT1YC3p1cODOBLkGgHB5sjrRsEV45kRScjZxjjJpcvQBUVL2/x8YCYYi9XHStks
/stWxLxs7gkMRl8bzyIk5BzaZc3aO4BE2eRJwZGh7LXxPV+4RKP0niWdrSejOYaj
RBO3VkCgjhOAJoTR3vqhAZog4UtKntOeoiVeaIKVoNNgbqeMDt5BD0u+rGoCFDBh
Solcx7T5WvKSGFKpTC5eAv+ZagonmLm+h9BhPcugnxcgz0PA75bFXLeJnFEQO/bv
msvPyeSTDQKoYBt8Dn1fpPHEALVRz/RP9d2X6cKAaUh9hjz+whLJqKBBEKgwfhdz
EYrA964s5XnERpTrujkrRwDATpw4N0zuYuU96A6x40HvsrMlTAVO0GYgCtVhC7CD
CkDU0LIvZYUwHv3CED/Xc212OcnN/SXHPRxMbLj2YzkA0iWh2irjLCiwQg+Su94J
QRl/p+wLR/Q520siPRDPZB0rvvtl0VqxWVXcgwQ/jQ95/YdKUHwjN4EYbrjvej79
LljqGDobUJwiAzOiiPDqlMZlj9sRLsTuB4ZONM1z18Kw5WHCntl/etFt9xTqMZ0x
bB9sX2nx0uvdzPcpP+H3i+P+JWQRUu5HKMU+MbpS6u38BZF3ejDbdjiz3p8uKwuH
4UHN+1w9AfHkUfC/h6ljUTA/x0dGipA31hwhQlcJmfB8rdYR51LSOTZZx5iyKprk
pT/FeKTTnh9RCQvbBNy3ztb2fCoAJ/9gB/tYGnWd4RX6kcaoapXueF9TfLbvOdbP
F4vbncU5xUTgVkyGX3qOHDpHWLzUWAk5LiUW6ImgsEf2TISFECWXDXnSLbkA0atj
DhjnpgC3XkEP4vjCx4AX+i7Od6aFexErP0V1Ibn0Cd2hqXpHdaneT9cSZJ2gVEAP
WcqvmWxI966RPR9jsOkw3Am+HNF/Tjq6PFznfu/njmeD3ditiyaVMHW1YSnd4iby
Ut0sPAWxJMSo9OJ7FsGA45zgVdDVjzm8vVjB8gTnhCQhgqK53YB+PhR9w1ydIJln
cNruiqN0K26lS2xw49iVydPAXjdWnZs22haaQNGUXuwTbTvacgIeMMYAFiOHLLNg
T4y93CLQSNPD+IRJq/OUAuF5RI0mfgbJQKTDS0dmbx+ZfkaSXa6uSoGurek0kzbO
HX/nff/v0yceYWkAp6SQpBuObPdhf4KcHy1cr9ho0cnIMfFXh2GHAnHZ9Kuzj9sJ
vIQpbT9WvYdn5HN7ZbRM4vkq/fFPrFzc10KKenMZbFyGez+gayREUF3LjQIPR0Bs
e6T0EUcWLDOW4oq0EPhuxIgi5CdtEE/sYb3R3ZvWam2ZpT7xmkJQGvZI8u9VVzXn
YpnU2ToKWuo38GUdyXBN3l6H9yKJgbmM8IdPiEBvdYTZ0dMJM23bwprymAlcFGCm
a5U9bTv4I5qz3bM+YLzJIEJ6jTBh559sDEGzlc6wTAS843PDHEkFQWAHsqdD/hjt
ilLB2MlIv/bcZ7t69qaAbY7AP8NoNSS8GsugO2DcZL1Ehpp4vdhsBIODWY68gBZM
PTVuFMlvXnXHZ/e8Cx4miQsxFS3he8Zz3S5wlB82ajjw6gtzkCejJc/Nn4FMzsak
Zm/kjl9h/5ekHb0tokwSdp0Xkod52c52wad+2mcAerSh2AcArogIBL+h69xFiFeK
Tpwsp8oDoSjHqlpY6hg6IiV6e0G2ZF8JhUl9VNHFZZklWI9zwiLawoCkWyewpDEG
6ylNWPVHaZ6U9srxe6h3uWJCawVsa9KpWWxqlnV3VQJIlE6syDGcARN8BzKZ40Bc
HOEOWiP0zO0MV3lHErLb0bofrQHbY1Uek4RkGm6c4AlCexiLKWcSQ6WEvAFPB795
AjqVqTaFFcDwaJJeZEpfpxV8OmRwwJNuC1lrtJtWjKYWpD4XHcYOSw1+z/TdgPhg
9PSO2rtkKJJKyhkDyXme7JwZDSZF5ETifZYHRJ6TTFvgur+1UjBdM9VM0UPGtvkU
nclXP/Qg9w1vu3vEULoS9i+GV9cj8m901sfX9ZQ4m8OIgswhvCenIrEJZOxyxA3C
ZB+5Rj406t3FJmeAPfmcGT63HfIBr5oBZ3y+ig5aC0nabuWKFy0ChMtt8iMGdyJ6
HTdSHQM6dBMusQ7vWpTws6XyCWahKutNksszGzNaFSs/YZV+Jey9C8m9VXZUOC2m
Fhen8KziV2/eS74bZZaCOfR6qV5SS860Yf+Yu/ag7aY/j49BkoqwV//fRod+p9AP
wunXmEbFqniJ/KjVnqQmDMn1byroic0kwSPMXXNtPc/yh1SVZqMYdruLnhJXKugE
FcSfoPmyz/nIR7elVuY0UtORLWpaIBoOhY/DFTvZQPcCvk4aB6z7r/pzNNwI5ybA
b0gPil3Igt2krivvByr2W5Z6AydzUEfKRalXieaYTOrFYT/kTSmAeC2AjhvD41RA
pjv+glShJyh0YlJVssp3e0tn5aazSM69EJvFaBAvwDb562Kicx3lbiv8b9Md1Cm1
4LQ2fAG4WIQ/LkWQ53pI4RTMSXgAvhUp1uZ8WxjXkft/bbfgM90lLPr2uEBHw9Ej
6zwfjPbyq6u37/UP943pIXqlfi4CsdetMIakKShDdv6CXnuQ5K+yX5LmgHDCDllp
t7gJZtmass+fpzOCTJR++jWZmG7iWm/eZ0+K1ga89U8p1qr6q0GtObW3h5X3eV8y
qIucLP1XcCqKPiQ14wEniknbEX9V1/OnpTC+xWNKxS2BrUSTjZXtu9TSmjLmFwtw
TOtDjCsgJZgf+/RqBLw36cC3szdqEe4BuyNZPHGm1OrBvTGuLy2zHY4nb8mrfFtg
6qFGAGFwFv/jJd0M7XcB26fNPrySvzTNJGKcmnVFTd25QVIBvxxCeXrBQoCFeGPr
VSw7KL1EQkVQyqdKohRfXWIUJucFRvB3ib8aOI+dPMbr2IWUX7u/1sixvpNR4Y44
VlsmDXSd8SVQ2oltWfD9/xvxJwOPr4r6rYVmuGO6P4A7MwG5fUtBgieDGtgP09Jx
U0IuxHAYSKLVCOWS/95kkZlyto/QFwTjSM4Ky8xAyuSYKf3yKg3iBBsw5mdeB1fB
xCUrFwbf0s70oX8DMYS9MvkFGOapyJ/7zL+JgwzVIUVreLT55hnWcWRbM4nug9uQ
6M8lfB/pN/F9NSObMKqLLGAS5SRee9nDOAbK24munk5cUfAjqvIJaCltBqooha2o
VunkdmLZQIB3rf8md0HQdXMOHwd40xzkUjN3HQw/MLvFkpmFl7dYJ5YL44ZKil3U
CSZpLbhFKm/c3pImm0f2VZoMcK4HNfXyFLnLc7NKsRK2Aagm+lQ3ElgwFq8eO3l/
qMiAppNlOf+6P+Qv8S5E24X0vMoLEHEKp1METLQdl6AV3jpA9QIDw+DDLzKu1iDT
rDQeAyCXD2DrFRHrriJZWRUZ7nh3Q7L9bgfCzroPr8E7Bh6PwU5m6GKk1kz8vgCe
wmBtvYJ6vZPjeGHICXeIHkaaMEwTS8gtRxuVOWMz8D5naYVGV6ZIsmlw5xtMtlCX
maLRcFcx5sNxTFmYgYjWhZPu9imgF9nt+dhclvWvl0FdFPkZAtIt04RWL1tPsYjd
tkAb+L/vE0nMfzOB0EHd5ExYjY5GTO6Xckqq1XuM4KAMwoJqb+4OzJgL0pFZNPgN
fv9I5hJ/G90m48r/a54uzUhtXVa50pVy0bepYJ82glaVVcnJtlPdjY8JH4/iIWte
qTx8pv8jk2NhxYXFdc+cAxuF5ygEStEARffZiuJ5mB4IJOf8MIZxxf94vsoNkA+K
F0duwIuU48soUS90ZWSIeS2OGndO4UnKMVo4LWZ5KCgPVCJLg+VbfXtnhqg5ljzE
spSZGKVROu0yVjD5O8RZ/wdBcTC1/OFyZby+qayTTqJY8XSkzVBCqzx9348tdIfX
YX2gpCFrU4Mrd0IT/clF2LysXVpo+i88koYuA5ios+jRr4bTQOmjvH1DcJgJ10jR
dVG47nznFesjMaoRU3lga31107f5jIjAr/yuhXzWFlLkVLc+XayF+3L4OE2I2Vcu
ocKUHMli+3CQSMDD4Vh0i0kTsTCppYH/bvu1zPDDaqjndljpDgnZlxNv7o+68GL2
G/Etg8DKwIfBGIr5FX6F+CVMSmFBBOwXHgMnHGgbDcOjF3HiON1joyLSCNsCWAV2
XtC9hIxZQft69GzuVeYkTWXpxgh8YhrrhjG9GwKhL3sFDj5cov3lNsdkzmlUB65a
yD7sZpbHbgkeMiCb/8o49T4H6aY8riAEYUE4pCHIKKw4HbTISkncY7fFJJ1k2vMh
bLuuDKp8eJVSPLmHd1TBhc4TN+I2YivuMJSK5wN5g68yhP/BeT+aaLVlTsZ8tXR3
MUGPizGbE9ExmIqFoGkh+JB8nNhQwWgO5HH61Kw8OdXOEWf0lpaMx/boOJJtLwzl
Pq4A0PBV8MN4IHGE7KYJohSwoX7k29YMoiOMWOAlvoKbDpuMFJKNcp0NrJnWADXV
YNfBZoxYSr15dzO9ZD3ggVdJTDnr9smZVAD9yv+JJ869xRygTTUwAgNRf6AptKUH
p5daStu8CG8eX/qO8jzZKXrtZMiZcRAIVoSyXCSztqp7iVVS9fB1O/5hcon7MFLu
lKgyjMFSmWMEB4wcTNySkWdC7si1Xbu5Ket0zOoGa35nCodmfQiAu726T6S9dl2O
inzfPwrVKrs7fz6sb+W7iXNioxdYmG9iY6l8VnFr63NRpVOe+M8zLiAsvA9Wnoc9
YyyRkGwxOBnBve2YrmboXf/0OMoFabQB5qF8sM84MYWsFemMGouj3ZTxAbfVQtsh
EDXw8UDIqC9FmOAFa5v31lkhKXXQpcsSeAeiEyfqhzQSKLa63FaumtjpvyCEvTY9
L4nTlLdUylW+XEI7zGU4WkIAKaXxFWdGqHtLe2XsFMnK1mmDMnc9AAJPvyo6hnEn
Uog3jwxWENSY4wX5ocPYKl2fTMnmb1slXkp9B0tEhFvIBCtSn4/nT++r3pJu+Vvp
aP9wWvJz0ATnfSm9WA28p7dDTRodQPj4MfosfULTM75hRd5LxnIix4J2+uZI08Dd
lqcwh603Nk4gaWlM0JDemf1TOcl1vKoz6dZitbSkq4GzssTzW/Jm1QQIvK5wRKAD
wtKwq2cpQ16ev/kfbzOGzZ35ln9MVS8P5GzpS6eXt8pDw7gJM4BUj6SWrb5TrjWj
9D4hHy2m8NtEvVoNYaWfDaJrykaHILuZJzdfIRljiWW/OubLWpUhzjYabdiJMRhO
GuMyY5osUee/A5g3bMQ8RKNdwlTE1U+3paG1HP/8iovjyi+NPGnAItUiaj9vvwjq
7Q+0ZZ2rBU648HMbAExSo80kJ45fRk3HsVsnRMcY2B0g92eH97SpQNEzlPYpcbGJ
orx47f9K47NbYkzMDoIZyBqtqNMqu/7NnRQY7EJAYEtEvEymGqu3R3FRZ5PMqI5b
85kP8xRkMGj7yrs0sA3NtsPFmk+jQth56A7InCfGEBmx7f2csOBH/X02+MzdtOD8
kz5iQmqDiEO7ADDfZzeV5Wf5S4zg17VvXv0+ynnXK4B5SsIGtOieB/+hRfURkANO
OXluiJ/9mH37wM7yx4uJmxSQ4w3gAAMuiHKil+6Hs0y/Kqg1JXFGDBthRTvdVsZG
Hp2ckYRfv1OjPQjtQCgqJgNyeYP004cKc/bO4Nw9Oy92ei7dsJHfK4OgjgJZZEOt
JYzKo+rOicbmXCtKWfyXJqqJgNtObGz1vNRRTHuoWvj4WpprrKqiLCVlja9b3MfS
Hxpnpm2zfkCsPbFuCin0zv1n63Vx00NjttqnK72D2B3B46jn4WvWP4Fro5GxKBCJ
38X5ZH0VbJjWquDL4U+mecfZWPYiLfs39RqktXeeP24KtJCY7epBHeWaLKI/lKdh
Kqjr5dESvtFOJL83Fu5rmQ/ihkm+GR7yUmaS180mMSukPAGWLNGBhq7HLk2s0Uuz
9OIBeXE9MqGvDouJdDrmCAJyc2JhGdy0abqfzxi27t6LSvfWli/5ZVt9w/vcq3o6
zkfkZUHASGw9CY3xu/VUMPybNTUJCwkKJzHcVY7+/EMg1Xc3cHXar0X0r1c2VDpk
zRcUmsCYG8wkSK5tBOuZeaRCNr/DHLsN/P56Ej/nPKmmiP0gw3WHAzQ31jS/eUYG
IbYtc1dRmAclQxXBmyTJhH0DjZAbq54Cl475qNoM+oaFv7k8Fojg6Atz4WCHVNuQ
/L3p58tCMO0wQcOKh63IkjndfAOYGeCNy7RyjilEGAJbHjVDOWdvFR0iZ8iBsxmD
QN3yIR98nZwDJ1X73V5umaJ+reeWhvll2lxplFVnfF00uhgbbRJIgsCEkiiEtwAI
BS10yi8PfKrTkJeaKvkkefCKATqI9KXt12O/uGb5wADj91mJiI0osZz3RvvsZJw8
cazoD+wYGotlt3+EEdoEdLOZiF+prQvPlB0MWtpkqvMp+idzxPvr8PgUJ/AhPwt1
m619HQVEfPzW7qR7xeAq6Hd3AHBLBQjxjs7S3Ag3L4AFZBP/mMd09fwcLEise+7j
hjB0HhLy7rXoSerT6lmJruWssShnvGPaSnGbSCEzag3k+t0iMP80ZXnCA/1BdvpS
HBiD2d2cRi62TASF7PaNlCOJ0CiV5g7hQmlhIx5pZfEoXeLQGsSah2Ixq0gRXSnV
oUoZikt2Ka6XjbbnaTduusJpRlwi4Ok/HyqkuohdE4PjwwOypdCG8FxGo3tnJ4i1
D2nPq7p+2Y74xgorWZbJnHm5DsGRdwXaLxSXJoVl9pnJdi6oOXYUfmGpg8KBI64D
VYqv+mX+l3areLnIxaY9ZNF/gcBA8XcJ5pKhoAoIZSG4/WPU5zhTqIimXJwXZNyT
2FcftcN1LzKUrjixnvfoDcSQQDEkrczPIT4+HE7d1Y5u1ls739jeB5YbJTVueO0b
lURsuMxWR7PQvVscReP6rH49VQZE0EY5ay0TUSe+I9L3JGsAkX1ZfszMxy2Kz3oo
xwVqnTMal8cohgP35DtFNpObhvpQLtK7mY/uz0u4ySyeYxXjooHFebNrrlHDCH31
UDA41N68tbZ9CrNWcYN+YSFk26EYynsB8XqF8nyWu/70auDnZ0X/q0x96RlxJSD9
wYtceJ8R3jzcQF6fHwS9BJ/+MqY1r9246ksIF7h1w082JQLv8ic59aF2OKfZIIMI
jm4tY5KRqlEzPGakU8tqQG6wHf+QW+pcwH4afaPdoIFnZAU1NyphcGyey9m0KU3C
PtoosvWDYxvulwukp85IIYLwZmFUVURlltncxA8bHm1levD2PWA0preS5veo9uJx
Adpzno8tPxHHUnlJoBm3M4Z5lYwuxss5nJQf4585Zgnm3oZC0MuZU5lXXHn5SyPx
fECEtM6kXcLk0b4HwStMblsBHyoSU079s1oyGVlzhIVP60/RqkXmIFvaJsWFvYje
Ab0O+dOTxpzC5KheErRJL1wT9QlJtSX5P8uZpZgzGOJqwiOCFCZW23mSTd6QbE9V
Y/fxIT+9ZnF9q0XIZJiECK/y6xCoEH6KZDzrGW3Ko4Mp6/3XiyPsiqNHnKLMIYiV
WTw/EZjqueszfet6LAC0EEtCfsImAW3QbdrrX8rTkSdPhucwDc0/Ucm5b2vgGZ8X
kGTObKBBiIqA9nOi9TaHz5W0gotKCzSEdENA95O5a3+4tInfNFQCRPfkTXVrp9k8
SSATeVccJ+pRxy7araTLA2/jyyahmETSJBaO9DRDi3HrbjUWJKsiAu+Bh5cye04x
6D4EwiB/DgvUsPLX9AOda5Gbvr6h80LMeundQbhePZaBhkihb9WulfnoNDYtY3tv
fe92i780I8u4ms2rdXImNqg5Ix4kdlSCXFjLk77qM8554gNHIqCWKQ7ZGnoDTm0k
iJqcPETS5ZGBOJWQdQoFHFwpPAkImeRtkQnmqvzqsPcEGuI1j/87BphVtbhB+Yif
O4h59sIryB7w4s5e7qiRmZM/hw8t2OvA61HZZqoJmOx2aMdO7xVATLQ8abfm3Ibl
wXAavwG59mGG44NpU2PjHYNlPJM/5W6UqJa61Jrh9Xwrii0VKPglrGTm43N+zGtH
JB0DiLZaoo1mADatIHDkfMtp4sYQJAvnz78gjq32Rg1KxKcmPlR20X16Auw1gyns
ivqouuwmy18VQPH1jph7Ur6iwJVj1NzYMIUshAWS2XqphD/k5bOGXgtxwmlQwnGi
tFU5nDjWzhL18s/Gl+LTOW+Ib2mbtiByD+m6pyrWmANp5IKynPMzVrrnP1l7LTUI
1U5VTIDej8wyCMMTYFIjUtBLToetF7d9ADssRi9IBMtbRy0Wx8ldnsSnKrN407E+
8zx5ha4C4PK2SGmaudvXjiAJx1OUE8X/J5YQNJm4AQyDStLjiBc3xXRcnt9k9vEf
CHkHKPnNk0K0Ot1TcjQZECZmBlNN0znWeTTYSfBKiiehLtkoc//EBol4zxQJ0ev5
GQW1FIaQh0n5INUGEMwi+I0a8hrMk0nHEr0TpVUryc189OGVUnytAi5O3mt2EdOk
vVG4XFLebGSg584NtW3+ue1hTjeiC/nVxi5RgM1cujV7YBbvonOFmTV7ap4ilN4V
PhsYj+MoSydLaGJpFm7PqDGy8a2jgeN+w0BZJvuk9CHTHIx9vGr1fWn/lmzqC/2A
+rPmRYVna/LR2E31P+j8Nqy2lWbCvgDl36x5lvmVYvOHWpz3/Ieh28bgAXDEhI4o
VnTXdk2qYNMiBw9PzDM5vd3WOdB0T2tZhzZHIrHeanPaVLeHnLv3Jl7PLASb4sje
bcUVkujAbVea7vU1jzDelkVTE25XuTA0u2wI1a2dhq8krIOQCGtbDdBYEtxDmkew
OxUZ7uhR0BR06K5UkZIgxFJYSY/MPyyQ17OlawntuFxxw7KwnbzeOzMfjgQqg5uf
2U8pvyfwoaPtQX1SsnqE9PmWDfybh6JH69fGaKF8u6oYP7HmHmW6niWqRGd71JGs
k3qjKFhQXrC0ECkLD1XwiGHskI4BWhGfOQwoBUavqCvpTrdIIWYwcIK4l/jxC0L6
F7+NLWgWWiGztD704k3Hv13m9xpcZLeBJ262jNxXiu2sZ1b2586KcUxQ7dTL61De
CG3fxRYU2EKxJ8xOuI3fekqhrGVNdbYcwOsBqBo74BDjJTTna7JnOhmZkb0E6yvX
0kQm6HkndjzSEepKi/cXCUIp0Fl+1fAaLzlZmh/exzIFFPArLCERrpkK264QOEnh
pygJQQPgCVgQiA+yq5G+Vtbh6bFisXjdZVllswPNYN4wZDkyuIFMQPKTSzZrwod/
InXqbcjcE7b7/k4XZaHZEoukN3c38ei+bepS1dyCNLc2sv2HSgeHdouJrg2vaoU6
LgcGGN79X5nSnE0ky7o4qqeDP9+WpnW8MC6lznSgY+V86vUmyJKprkwFhSwVweXe
IOW/9en8JLZbBCtfmBXRd/VD13jDtdrqscK13FwbF+cQReQ6IhjYcMDSn7DHSLD7
KAd2dR0gZjQsdP3MZxWEDLjz6Gk2MrwVt9I0+w3NGl7wgaNK+mkhdTHdFaIvY2km
/k9Zf5yVa8e1DsiBU67CTat2Js3+/mgcNa7zdtHobcUNqMM1pbsr1ZEGkc0UR23c
94tlzLQppfPv+QlxcrKHYx2mM0TgzCyhXSClyBpzDJylrxyucbc1wKaYHytmb1Px
MeVypyzK8WicHG4yKhT76pBKegti6K6TGWQt9SW2QEtKaziey6I0yTu3cpVO5FH3
geKq6PhFwqlNOWBGvxwmaLUGOvEiCQd+qroocjM2W64aJ5zmbYYnhTtn/68nBB9B
hMo6ZGwmo2Bn1s7liiJ4YxoCID1Be5u5wHY6RoXEpCXPcZ/9Ms5ht/TOoMQTOlGu
39lAFI5TDkHqzsBqbdcL/gBkJTYRSwUFpRWhWA6Dw1csDHlY05ooLX9kN991wafp
tFpAnjMLVhZnVzXwdthL9lKqNf5QItIqqFiAY2+5sDyMKaxeditv5IqziUGUT7E2
PmaRkfz8X+aXC1yVjdKKThMdKGZXH6Z5ennuNGiaAosDYMHoKJq6dYwypCrNhgkC
s32xd1S55X+yibUqgnudB8Y9P57tn6Ptzmo4i91f8nQKv+YB/k7Yg5ZFMeFRBiu2
r1IDiNg3LXTVKAl1egEU8GJdIQqdEmsn4xF/DxuTVccRf94oSWL0XYYf5mcEcGuz
TsIzsirZSHeAPeeLdkFBbe1igGqsea1MNVRG0O9m4ZwQbWqjVIkUBvJX1/pgK7Xx
Y3qTN5IFZZMVwl4yrCG9G57U5POm4vRIaBDqj9GzmWEB75i0nytt3kanG2ihntuj
bOxg3dqTELJoTjsf/U8IHZuE7T9IjRqW2n8UycBFCEbWWVaXiZ/vY0aKKtING+Kj
ydbcL4lDJWhg3KlLNElWYdSOi1DZ77eBMBO+FPzdjiYWkm3YwUzuANLJUTBT1jZd
9TcNnx5HDRLq8onNRsJLrhmtXqRq7ke1vWLjV7EhA2EyzCJ7q2NSsKsAr2hyQIBF
JkA0L64K7npaLTW94MQXxjB2KyHSi6g4Xgiq57ee+oyOhhzzBg+gWj0wDSwgAcsm
DnRjjpL17tYy/wlhZYlHaeU3R9nxab8qJz8CPQL2oEpnIJ2wRMmIQrUm8Xw5Xgef
4RuJ9TZvwFGCJqrdpIf23KhVzHMiexYAZQnYZgo9zf02iY16RzdK8m7hQOcFzCOh
iio0RZdcTzUybvYr1pfy1VFVzwiagTOL84+962jsauF+benIAUMHQUMw5Z9Qtbzh
r/hbdzk75y0PDM0uxZrnGltNaBn83RTFIbRC/6Meab3P+6ls66QVtNFI2ChJyQ2R
zCq8toLgOGZqA1glk9tNeehgPN7KNrf7RjUQ3JWCfd4FtS4/i7QZidSnDh+4zjzo
FYGIV9m+yvRpsYxw7ETlueqFdEBX5P4LL3wk2qk8jM+B7eCcwGIBrwX0TCPjy1c7
VNJUJnIyUX//xe/2/k6qzIPb+/f01fl3IoVhSx1YEqgP9fiD3nSNSYy9WWlEglod
zAS2oNOwbEdzZhLXetLz1JICVt32Z0H53NPrxKQnuZSv24ibDW4BKLRz/uHqR6iK
AxqKGjWRAPOezsxRcloBDZ620sfJKTQZa/I3cWaup77tA/Hsu8/jJ8cZF/I3flPk
kVFN1p/HfhYEzrSKcw08CUyiHZL0PVHDdoCWwkyRsOE2pKYCaL1c/3er3LIzv2G8
G/nOGqf0Roa+/1F7vr/T0xEyFmvxbWuGxevwJP2usL+aS3ZTYWustkvTBCEKRB0D
csDCAWAcDUIGxV6Eml+HMwuGW9dJF3ybQYBU1duoeqezCays+3wqyTidcVw4yuL/
LAp4AqC5qaSiW1AnNofKxefY3bbp7KuGJzZ33+xjk8CC0juRK6avkUy54zSVq84D
/Q1AWhR+bSF6XS6g5wRdRTxe/ot07nZQfHx92C+dbZvFkiBI5X/r2Ws3+6qdJKKv
6RNan/W+8gXCu8f4oE1DnfRyoc+Dg9lf04R+YoxqNO5LUZGD9ogRVeHYMNgswFn6
c8k3nwrSHpxPFLnnPB9C1VN679FLHAuDNXYC/MHNdIKXQsQafijq27/lRxJSHn/G
LiwVWXWvAHsz4m/4u1jJIUJI7H5JWZJY2raPEINBOhZLAeMmhT+OSXgppVczNXGx
z3S92XW37OycJvXenyRymEIk93Z1bXzINBE7kXK8L9gPbFQIraCFc5RRuWA8P2P0
lY3PVvVckMCPHkM5YdSyz+433bU/TgOsvhGMDxDWuY9fc/QN2u/FTY5mGltwo2h+
TxLhnv62VlSV5MtkO0h5uJHx6UzaVXB1SU0Ppm8XcdF6GKZRU3RaGi6PfTX2UT20
8WvYISvv2oCpo9VXWix48kiinGfanKMHnhDQRgvWpLEl50xcK0CDN21G/SURLn6h
UH8/P/jovvxzQjI1yhkDYJIcoMnc4FHB/bzZh2EZlr7SuziHtIV3UeJxo02tuAGh
WYmMB34w9jeBBigd6vsa8/qU0D7etzY+qbwW+9M4sW8GMgYuVGosW1oxkc3wUodp
rsNysXXV23MTjTujRa+wjQmcFMjJyYq9Ta3969kQDC/KqA+DnwxjXHAHd0cHqEQ1
u3D3xxMBu6N19yXUJHEXjaYtPKpoQPls8AEDxksQdiNcKyzA0NXnv3NKynWP5m0n
F9EPWTfQoGHNDygjKdUMzRXKaE0ByS4gI7Tgvo7i5gvsQbgcox3qU5qpt9cSO39j
7MXJQ3DQqRB/YFdQxBj+mNTSabHJ++NeAxL6BCqSqV4GH9LAjogWUC+liTRW98jo
7WjC+fwwoV5g0jLW9gt/zztPgYHGKUbFPWlJhxCD2utJAyUTEaPxz02aeZGDppJa
YwKvWNWP8CnoA6NLaLxXzIGaw7C+rA++rLdQS95JvqD41PzInrSa9PaHBL/ukp30
UeWDoz3ezM/ABHTWCRebkTlTXY/5GPLKz2TfdUZ3LFjPejeTBGSyHL43bEPfuexZ
SCvC6vqPyZeYK9hInaahw4C6URO2CpenNHy/WgEZ4DqdgnMD/81u9E2IVuuMJt3V
SXIzcZcNpUv+gMgraiKEu36dEryMykTzfMHXnBaFqGc7D+9//xAVnEVmiYop/Svp
VHI8MBFlfSJd8U5tnmjQ76it/ll1Q2SOPF7y71rBTtVDhUH2afXF86RbPMC73aNB
wpJAisRtQCcv/yDOHwqU2QSNYwX1DiQD4eLVVY7rFeCDP0GYX3sVux1bBPMqK2s2
9dXYSeqNoz6L6ZzkxFwWwSLrkPJocuYwVeiHqMzJNhRVBFc0tNyjR67eEoEkTLQI
z0HF+AT0IZSfV05w3eOaa3q2hEPmnlR5MNn4pGu++B5Zs98HufsBWVM1DpJCdl8D
d14I8OAOguajl5COBBhlRYubSbbt/MTxJtlxq8+IWDBFHC3xqebWaotHmG4bZzfF
FvT/sqKQuWRAveqeQKku8TWw68HW8HegOcT5BmmN3fObsFwThXE8YSHbrhLoHnT0
dWoytb0ACz5xbhZNmwSbifPoAZpLow+ECB26A6E7uYqZpNl24YHLBTeVj36po55q
peEc/h9WxH8LzJ9e7brk8PAV/cY8bmzfQFTnataD4Wj04hkDdPBuK1Q29QmyKHU6
4alPf38vYnoEqonzHHOQIWfd+Pk3x9zJxfWSWAPj8WlN4CMesX+g03jLjuiw/lBp
I4eF1bkaaqA/t4qFQ1rq3ewqF4DRjmGArk+p8N3vhTkiJGtdExVi+oeiukIB6Js5
oaZgFjy1qHb0SxhN93dIIgzRJx+XlciZv9hUUgA//yg5/mArLoRw/7xjnXuDaNe4
t+Yigz+ztYVpTaO4LRTa9nmucnSIO1VnyxxCANxCC3vJn5nX09eNGTUyRGIwdnKf
cHPgpDoGLqlYsP5elzBMN50a/rkShfeY7tACZBIxMfE1Yavm1PMHZXM2Hj02/fW6
y5IXqg4uttcwWEHzarTdR2+0ZlDtTAlApYVaDOPG+l6WRYFQ+uNFIHPlsgn5EFrN
BKmD3pOzTfj8lPAk3a9DNCZo+R+7e/d1vLPiI1snVwDmKekEiZNV0tcRUA56ERj9
N2dQeXbt5V+JPAtmOl4mSrYxEV8KhXMW5m6x0fjqGGacQFHwXPUk/SWYgXn14zrX
mYX98r4Ez8+wUwqfOfkf//+Hgx6IJjay+MYe26nz7Hb/crQzc+TVuRuMfaiiPyGz
o83H5M8gyjCnd3GHLM5OTyFJIReAHpm4J1JyBBu9v7VW4Q/E/2+oqSvWTQbzSdnP
fAWgtV5Q4XYk+nVZAN6anjAFQt5gI+L4Dsym/Xv4Je5nIaU7OSjEzunTukVmqTMW
OqlKIGSIFpPv7sFBwVH/Ogbr2B6sSmQISN7ytlTbAu7/DKnGDn4d7fqfOR60T6if
exI4LZuxzFAysRLIdQebWSDFjR+OpsbI3ViDSdYx2Juu6kgPD8H3ZdlN6rhNmnDL
/D2g3BUleMV1d19TxV/HD258N29QfBlCiciWK2rc95aEjPI4hx85I3NOgS64xhuI
2qBAxk5j/r3UYXh+t9quXdWMvAUYvxvuWZnCGKNk2fnBuagxuXotkRuRF3J6+t1u
rwzJPqCHAVEYi0u/GEOHHmKAVz/hfyaA1zdOfw/UCyblW6kt5ReLgQYdcre77lBq
skfYC8L3XJTQCgkLIPRMHNlumHSHw/2gom3fOn23xK7wyxfbN35bymTxkmqAhQhY
sNRZBAMXkMISPwiaOuE6oS9XqDPr23QzooexcRplanMe/Wl5pTZM712Pnrhulm9m
VJuTPhvmiqkKYdmffjtUJhu0OvBrgpayw1Q9ZncPt8igo/kFKu0ax8mO/zaGmBiq
VneYKbsthg3Pw1HEtJCqlYeJIj+YEHf5Ep27w3KI5jZyuSblAOyUW+IhsgP1N7Ai
7RzXerrMHB2L2xc+m9DBuJqhwt13uvLW3o3diN2P+RxZP5sm7jgmr4x8i4lYHiXP
M9Ocw82IDR8+hb+oUjQGQAC/Q9wEsLFMw9xWWKYsVOQ1yHRDsqzvbPONLT89qnAK
r3HDY/ccyide89QuB8EP2NN03iaex+KJ7dXCvS+3HVwJq8NpsRXL6XvzP4s4/+rx
6j4kvAYou7lUHfQ1m3RO79jeBOICfDXULxuY6lMALUhfRBdWmnGpTw+ptgHk191D
6eQUViv3awNSndquSITSdnIwBwcdIdf62VyRsCdj2HjtiJPWpnPERpBv0AwmEh/c
FUNbgr3J1lg2ryYIu2kHGkx0KSwKKkEzxJ2uhzmNy5waPh/p0lsP1/KL48yo84KI
zAixX3+OMhnI90pNRkdecrBAu8DLb69vh2aBsNWRDq8c/tXoQap/jr7YQjLe/mZT
T9YR+rdguqWU1QreP0jmG3B/1K5+SKIzGoKobDWsAI05fbFJzvLtU6TfygvAtFOR
CtQDV/WRQllMVRlAHzBeqsjy4Rj/R8jJjOiMk9RC8kk4naCS906HIJH+e4Q+qeYc
ubc4i0nCLSGV8tG5ObPLVA2KBqb/nCGUSAJQ5evDXU/nh+FsrcH/cpxBpXkumUhT
yfjWB/qebFPrlzJ3XQQGsu1XyVb2nxRY5m3Se+T6fLB6GxBPv2mzReoz198pARsl
Qtg+vEqHtW4hoYo7rwanHhq2tqEQgvLa8Bi3J76q5TJsJZGIgmgIfA6GibUumOW2
fL1KwV1pUavZA6JVjZnSCvEdcw34Whmy1J0w/YWsc27vdtlHfT1/gxcbmpib1GS2
Zq693vaYnvFCH5pthjVi/JNYY6FT5352LQWcSWD+UnLNABfVQAu7a2DwMZeA3Ooi
EYiLpwhIi3W6om0wSeaUWKnF6b410KqfEDofQG6v5MrplreaO2BmDrQlvoAb7Yvz
1abcTIqu5RWCAa03HFcqPGZDtvuDZaWRN0td+wYCA0rX8INLUhZOQl126Hgev8kv
TNlppMN3YsXHl3E0iXfABv4p1IUiLzXci9e0CQASIuNWukZxqzXnFVtY2ui7ayU3
L7BEDibq0ClJhXrnY1ywqPW449rir3ANryIJzldwo/RpC9DGAyILeoJ0TR6jmqYl
5A1M0sYIw2zE2MKvlvbFyCkUg5d3qNpQ7NZuQ7PfeGRtynvLWMp6ski5m9BP1U/f
Hu9D9lPo3thxv5P6o4vyhZzTUn5uKGmIaSsnfDx8Cc7VOFzOoFr4ZXmPIRHHrslr
/vQCn1qWFYNmNnG5pn0JlY4Il5nI7YTcf6CTMtknGDHTWInJeXM9yILMGWEbGVz5
QgOyBWb7Ne3gytXZOhyfWYrQUsX9Mizqk4chBBYpwi5bEm7kOyByhcJvTvtjOyiG
Z9zudVGMEU3hRkROxMrPwsNYFuJtcGIE67xcSnrZUImz6KQFCwl5aoY3NpopX2pl
2xS5M8UY08tl+qM+G9BPFxW1Meq1ZI28aPbMtFaA7LEqIRL4C29L39C0Y7mo4mw8
BM3rAeoB4hemKjDuIaKmBmZJAM4KdSuBRJUg0Fl4qp5+8knA+0zZJtdVqBgoghP0
0dfZ2KgYfN6s6ww+ttef/uKaqHUjePvHtd7q9IThbAlM1UW15J+C44GojILBb+wI
psXuaUzp6R71arpnQOeoNJFKFJ/8vCMt8wO0e96IEFC/P4K81OPvmzjxYfw0axFC
zHJO3jmcA4zZ2C2E67RqBr8cEo7qSWDilUrEmbjlHyqu3pZzp1z84nZeXhRUkEv5
v/tKvOzb/rBbt5SlijMA9ewnDByhhONKBQgTyxfdLxlbWwooSB3GaubZ8jhlnf9K
SXhySteZI28W7CRXZsOVDAxNLWmFZbM3IpU8yMJLLw+QEKDVXfHAgh2GbCRgx3HG
qvACHhwI5YuKglqIefk2rboKM2lA/GTx4MnL6bMIAGQRtjmSWVJA6wzyDFdlRS+M
Fxhec9EWQ+g14rl03gMmc7Qrkbdi5TXLMJR9519NKjYb9tR8ZSVDZLV5KccpuLHM
17pQqKXWf6Ev1nTxS8Iz1RFkma0L2kcDt0peGCXwWZia1Jlp1jXsXJLNfY+Dkr3S
QjqaHEIitlF/QMWZMOFQ5qftfcmmbwwk8zzFXod/cIhOuXFGxKR66x5NQXdYYMru
kJ1E7wFhPfjuT/PN0X/+4UuJ54FdOs5t0u3Wo+c2iWpYLK5EImPOmCEQCNZ6AkO0
/X10rkx1HwZxNR7mhhpMZTMftSuXzjKAm7M/fuxl0SKQcZ5T16wvIz1T/Ljc3kHK
/Rh+D0t+fU04/NWAIiCwaxFgjL2FxGgrBCclFIH8r+a+Li2cvRZdISHJeYDVUT8W
JmvwIAMLl7+8pKxZxmUgZ/M0GmL6EUwTqFl0ElOyvWTA0Cdbyl6wUIre2oaBt/Q7
VfaafcnxRV5+IxbKEfGZo4NmPbRPVs1VhpZNuOKoAZCuUkjNsZ/hQz4XjZ2i/Rhr
yySFYIamSvKAn0l3biY+HBAFRvvlBgHkAThPL2up7Pn9UhijiSsY0nsJD9dV4Qk/
ol599y4BltTmgq6tdjKWreodjtAU8ShOxoaJMp8Cz9W4glcIH6yEo8xkNoeNgve/
LHQi4418y1qvI+ToGxUsS+j329J+urbEJz5A+GUobiyfdK5rcGz5rieuPr5v2xfm
izUyKAWgaLUhI8VJhGinY4zvVPLLz7MfOukiM+jXJFsCeTZmO6AF9KCK3MAnhxNq
Q36hajYNlp/ihWj5NWqiDdzoYT2KHra6GeqVF3Pw7Od2pUf0Y81FcGu0bsjlZ/n5
dZ/ZQ4Thuxb8OQqtWE3/NqYwIDkKF5sCkWy9SStGsp5oszAJXds2B+IXqazsomvw
Z8qlH1IJUFqEqy0gchHkd3SIXg5jI15Nm1Q+Nd3uUdB4X3+lAuhmj3vahgZ8E8Re
vaFap6cZT55ocCGd4r6wiutvLDzTWW0v1hnW+nffmy5EPqNMGfojnqRRvd0x6dCn
0SePFO1oAuHmQKyqxVaSu1BxnqV17+VzFCSBF3OMSGVVoZAr04Pvl4+V2ZevvAnJ
T83R0/0ktI5ZKv/BQYo01FNB8OJgABkHheDPH3/GM8ibSP1q4q3WoErsTzMfQH8A
D+jWDCP6KdRVvDcHMdMbH45ZSsbgczScEACiOJdDnpuUg53bxkGOIf4FlY8Puvds
dJjRviQtF4iQy/TsjmVa1lUMSKqcOYKHbX7o6kIjEQpEUDQxLr+jCF7vTu9/4dkE
jVqwSXmUeSu3DHBTfrpk+zkDJL4AReNw5WxUeo/kbQ7wXzsl6d8uul9oWZ4q9gVZ
vIvNP9CduqPWpCCh+ovIJqQVra+JSQsSygFM+rSlYQ3LqZ2lQMh2MQpeuwjA+Q8/
Z6sE/SzjMRfOpU1HUzxu9vIpejMvWUULkPSFeu4cwZKm2ZwEhlPDtaA03ygl74WT
e45BmDhIhZwicYbTGeSIqSOg1UHPixgCBYee3WaFHwHTbbwvf7GJCJ9y1guY9CTc
lMiP84qs5C9RPpjCZNLhjG0igxRf2Na7O9X1Wrh3jRoz/Htiwjvngb6gLmbtR3De
/9dsskO0thySmXxWILveDYFMzqXx8it9MEIxmT+io3cyqwIwlMS2AAfNOmpi56ug
bF1pZ5vCm5bvo5iGVlpJyPex6wOV5FlTLi+6uxV27B8koCLe+/gjfZtlLdq3hojk
PmqYRBCcvUui2/TiHLx65fNdqydpgylRthEyZgmxZ/I2/nu9FOlrzSy/1vDw3d2t
xl0F8qzEqnaox1QVvTqeTWUgVsdq+KF2k6oaobTo0ItmXpp59LbdXZDdIYAur8Zy
OGrsh6xE+HOvXMgLhDoNb5xfW50baaAjXa3pZuV+fprykNBiLRqFgji3Lb2kwVzq
UrUfzBCJAj+Z+dQ5NZSkyJvkcExIc/3BtNlcQaSXZGsHMxIqn4NLcrKAbdYuG89H
CNZVKXQhxYfQ1YFx6eFbXg7gLKBatWIBsv58ZpUXhFCl4duPMP5mkTwi6P24VLxC
X4rxAB2JRlNW0tKRQhXKwehvLgQAMwB1dY3qbzCIiX5lcpwu5KqaTUDh0I3JoAGX
/UQQ3uL0PhPxtdZ3D8dkbql918vVpRJvs9sKE+KPckSIH2q5N7Rr/n9EdCuWsTWF
ms4yndzmZau7/tkr0aZA74QcSQesLwmdEeZ9fNg8dt6vMUCuN0HogGzFPPapUvPw
rU+FAIX0vgK/flN3ArPK0MBd02yf270qbO8Q1DvnlnVqI+EhtGUXk9+Ynz1cW/YQ
t0FSEovw8svwIlAz3U5pDqngNAoMUpLry2eFe+nbRvf2GsJpvisDBQrlkpqj4CUc
sUoUPJ4UktH/wxUbq9oAMCwAUyyXnwJeRe3lmOV5WJSeHzLusxK2kHVM2IcAC5l+
3pUBjuVNaiWKWqssZenpLwN6D+ZkNqKqEf9B3Vq9ah1hvEnmPlOGDzIq5eHashjr
ffgNkBTB9bLG2RilkD6+THFp9td3JDy1M/PDXmqIVreuwM9vjFrP1+kKH8E6hohW
Yt5Gnw07MrMv4oyNgIIJrUKdJFUOxR/Jx1mGUw4LNULTCfqaWyqUtdKBNVzy5xfT
rssCyBQtvETV/K2S8UJOaeD89e1P+kVSPIBqAA5sH+B/NT4Bj9TnHpxPWZSk6oAK
6MQ7xu1ZqRWmLDHxz3HXksMY+L1zXsZtxRBT1hjirPIaHREYOo6lX3xLkdh3oXxD
ckx4bUEzw4GdLwlg4etevhwRxjCqKtF4gsEUa7+nZp6GvOqHsyUINRGEGez4LRbO
WX5AQKPjLlyxrdPsRMdIxl9KfyqTJXmDnEBb8kVuXfglS0u0VVmweFftC+dFJK9a
p771BxHE5B081bu26vyYA0G5QxGeenN70JIpGMfrAJAX+0epPRF7P4W9dXdLz2Gv
HWWCRN4/iCZ66TcRUC/kSlSW3dGJQltitTNT+r1ivzlmpVCLYizGVafg4UYcQLkJ
237Y6LJI8XqW2doq830Hq+Em0BA6l2GdpOF2rNW3+XBz1uk8WRBjya+3neQedYbk
FV6mGMZ/aWarGevGwO/Su/HCiUCIMzfgFWdTyVM1Yv18JxoaXH0EsvWZUy06RsUA
KpYDfMWZE5nvxZ6iOtOFB9ZGd9JamoizlAs16cjeXiA8dfJuXKWE9K+tOkRPxk66
HQTry8lEiEmOcGJIdAVykmkgU8mDp9XZoKwy5ugL3GH7mxQwI6HAvpfXgY2MFqwZ
ubyVkjjcqCCF1GyIenDdjEqzH8ZECHKd61d0mkR44f5331BFo1eE8uIM0Ex2/a9Q
yZFDdpX04n99ZJPaZZpt8M3xJAoTJemwo/+6zk9rOEQwOEh2F2vlhshF4dcE3xeh
N5ewfQzGlz2v7jbJMe0unkxUBsGA/aSySSXWzDQ3B5KMEGpVMxaYDDKt4E/BJzc6
HUGm5VAEuGydaEx/DvoHWhIlMKXgi4h3gH8Nj5e9reyqvzfUwdUKoljprEGoYoMM
D5h6k/3gKn3Wc0OQbv+NdGgGkXwrNpz/elVZhGtaEbsNaYcI+6wBjVnR/9pVnJ28
pxzWY28EnwuaK2c/kBnCnYw54Aj2u7RR84VAgTm3w+zxHuD2lnJ/p+DNsfQVI0Cf
6kDwV95knVvexz7dD7M25kgCShZF4H5PPFsayDsEOQ9rH2B0trsMo2uQ+oB+Ox0L
dvsOvRTdfPGLClAYFb3ievLsQENG8r8UqeRLB/MokZ5qAZIE7RFR8U61nyZEHxpJ
hhtr7EoEvLmXXJpKAIuwdtdvG7jRomVPDHrK2OIjeHlSA7NllPirsyxKZjHa4Wwy
5Ooyy9qqe/BAEIHqVS1ZBVqx8r0tXbTubrXo1Q0hrz0ohRMk/aKfLM29faF9U88x
wehzj5yFSTqYxcwJTu+TVKQlzJnfDOq8Ei2xtqdL561wSom5hs2ONBV1OPFP+nPU
QZqKCgWJL5oJmth3LcQxVfHLcdn0/JbhrZgXui761Q7Bv/DJW57T6KPVJvjX7Pzk
c+gwVtm/Xlkc1lcBiTVeBAM+1WUxm/nOeBFYj8/7KnzFo/JOV+ktqSWZTPEq1XMa
nh0dLPnJf+6d1qRnC2Rk7P06Y8Fl8GojapPEH1Ppu33ykKPVKjalDbwImBy2LhrM
NuSdZICGWY+vawACe6iO1ZTA4fzq1sq1GCq+tgxWwmMCxp8HZ3fAETFwsgi3WDRA
7mANOOP3nvRhQP+09gVqM6ADjKgMMN/FbUfqkv50Cw7QEuxyLCDXmPy2CLCplSLV
MLhmztWGfD9CjqOdEspJ4d1Y3XSbwK809wJC+uviTwId/zJPi8+3cw5Y6ccMsplK
M3NzsfgdopGQmenW/8qqkHd0RM4oMmkytLfpLQBSOvMkIP2KJVOAAb1xjtr7SN4R
CR2xD/LwPLf3ssZwCsICQRzk67lOwe504WTp0vN+PzHHggxq7tkBXUVKJWz7QGgb
ZnkJw3FkndoLlw+5ic3BgEJbVmdt42QH2SAN1FE2rthSnMVPecf6rccxC47PuLFC
gDciXu2S9THzFLOs9bC56TcNLx0RNChB0w0WpRHvwrrD2pvQzLoDmd/tOyLaDzs4
DUlcX9BcCIk6xFj9PG9s5fDl2F1pesmqq5EfmDYqX2nL2KSCI4jUKBWrl7HjagRG
HBtjAco+BuIIwwl0CyZsgXnoP2i4RnPpmzsFdD2q2SwdRqHMRvXueAP2bPTjJLSm
D91eoHyQgUrWQIHTF/4tKL5lbuR5J9k1zx/BXkATzy/9FGEIwvztoDL9v3Wrsi4X
r0Rm1qgZLIVAUSnLiInPZdNAmtl8OR68J3bQKX/y5yTYDxjr0tX7VbQv0ET/uTx+
tNzjp1uTglwUnfNQ5b2+7xj2ksxC/Q2/9GSO7M0P2Ewb0ojgVEFhv7jlNs5Zq+xP
jjAd/W4RUixol65flPEWW6FsEckel7ZJaMKZ183OvAXzefGiITSgnhwuBt5H9RTx
++29IA+t4O5+QE27Q92ZHe9Rl2wS2v/3iZuafNqmni14j3/sXrCrA8dpNmo+NDj+
FJZwnTOj93nRq1bHnx8ukhubiwBDI1BaVH61eVdHhChpjWUwEMei+Cqxp48KZ7nv
h0VryvYnqTPEuCIPUYVyle+4shxx4YFyJ99v0rkqYjV9iWEkT493OZZNoHVTbhvF
uM447k1iY02a8TLhOt59dYkIthIkWBtfxQrOuYATe6FRQEWFkQ5LuPBgPalqP97h
rqJr3ae8kITyq/tPjFHi44x/IWnmigChzXmkUiMFwmcRGirSuV1xplI3s9eJe6CJ
PuajQ55fNoY6snBYhL8ZwDl4F/VIvZ6I6mwH1Trt/DxYIRl/3+GGtc750+dY08HP
d1Bebf27juIVrV1DHPO6jYpqgsBa3tcwH22o3wmNb3ShYD/5pA71T8/pfHKhpdV1
5Hl+AJ3yzwGwxwZa0YEbgUm6DEkRGUdMN6LN5FH3CyphEOb0GfRYUoLAXA7rwUHi
0jc9gS8qEXF4RYx1H7nOyQTK7X4vREGZVCLpJO8V419NfG2ir6+FWDZmOmpR59qm
s1LnOUnBdDkKJr9qqe8dnHgXb2MWlDbRcYQYElquBLWWI5ANdQjLOMzfEZL5gOgY
K5bIliBW9SfvhfOmXInatuTP7/XZgl5fVo0nvuD0w3gqxzRbkWxGO1W3dvnHT9Fj
8W3hcIz1g5241Fjwm2AvPvkx1eoQfAii0Hy0RnQdVtwKhlCFrlMQ4CMwoIUTsLAz
Sr2V1NA+T1OgVc70v0LyNEg80LLxF62CSJeGBh5g+IO2krrYOjdexsJ2KqrYWwvk
rXvtALVe7Hjgl6GGWO9VtsN0abd1zmk5yZRNpLKxRiR67Yu/LedGQKTjdE9sxdj0
I9U2RZ2vmxqAt1gi9H6ByDw7TQ9oc2QTRPG2FtY7tKaa+Nbkqdcy/AaGufNT+n9L
nJRi1Updpb4jNdvFidJU590XffpI02Zavnb/R98H24p+qyz/Sj5lBonwTnhlhtn3
bnj4RNJfw1GYBmNr+Cb+D4aID4ekME3hZ27NWvp2vwqDsU2y23g19jWu8/Qrqhpd
muP+gdHktDFsHGGMN1wXEaevOmPgAfQ0msju0Ax1aQz6LayzMloN9wCAiVsOYCBQ
ECAiuSLkURw/e1YgXH8XaGWxakrRk/qRNfFrVGIU1zJTLYegzATr7QIHdaBLaRIY
9IzKyC7A0SoXgagV4qcmhgPaxb29AsXpKJ60kKOsNzC2f2C6Wz40voJ26g69K0yR
8vvNvESL+LNSpl82dcG6uaTpLLq9Y9Lq8Una6xKrFA79wHD9WXxqiLjtNnaemQD8
SxM+k7zJ3KoRgFfqcrB7Vsy973duv/lR96lMkuWluKsCSbIAY/2E9IAWssD4slHH
/s/SRckDBI8jqN3Y+ZQEvlp7GWnLbxbLjsyOEAoPXJBzKHF/Rdc9rEQQ1VZsIrn0
JXqDdhvwqrIundtXi5NI3uqyyQ6fYicnh0biuYqorJ0iEBclOd9pj5wzGMM7pcVG
dzO2CagBTlkjjFQM8Z9RJW3s8KlMTePpgRpO45fz/tyNFBUri+GPN69W74uzGmfn
JrrepZLXjqTJiuKst4C8aNR+6Xg2Xkyx0snvJK1sKRf7/uSByASkxuIJLDxbJbGL
TMX+putYzTxmK5VMgUiuF2pbL32wEFzzUqFFcGcNulhmpFG/7o2wvB6SHw/KNYx6
kdUe/nbmF82ScEET8dFEXg8wQNUKV3VpUSKqyoAOhg9JPT9iIGMZhf2fPsSc6EVV
SeO3oYnn+VM+tx1Z085MXA2teIP6wHz6RL26VsnANn98lSS95Vr3+SEkM/UeZ2/n
jWVktsRDBD6Yt/Wk80mwFucwcN5r8sy2YUVWJcq6HFLUlz4KiDvCHJUbsT509s6H
aIPmefvp442A7aKksHKeG+VMbtAMiOb3MjYKg60qifMbW2SSvu1iPvvY4E5+Wynz
5X9X3gq6FASpn62XlYp5rewEzbWIXdo5X0RixdkHMaNoO33S4HNX4tkX9WL0LziT
3kYGQ6GhAVr63X8ReSRacVdzcpC/GnUHEdCs3EE+Q0c3G1747FjUS3UyWmjLodxC
FQNur0pOgSNTQrV48iqjLc9tq6nlbjtLVRS2uqxE1LjlnmAumueW+RblXr5NkKuU
dxzttt8vf3hXYE/k3qqT8IaWK9o1E55Qht1Aiqy7oG/9aRYo3goKDTXsQNYLwPZG
jBHlQyfX47MRrwyWy09Z4RJB1cQoV+wPBWX38po7MCLtMqfY90eYd1+wFY2sT8fQ
NigSmXYEPLi6l3mCkuRPs7VEAW3H/VmOQIaDWgOtsFtwh+Q6TSlFdkhL14+Lfp0h
Q6EXBQq2vHeQJfTezaoHXzGPUte/pc8l4E3RYlV8V9D61OHMgik0JbcfhKVm6p3x
vBhwb8b5lq9Byoyl4xbIc2mxip70VGMOfLc6spLmdeRGYxqeiZrleUIvsoAYSMe4
Dl/VfTETYeC+2ctdCCjM9yVU0OWUe1Da2LPOyyI7jW7NdL14kJkMX0Rz2Btg5Pg3
nv0DHfzveskV3A7JW4kY87tHyCGIdK6LQ0AtIuqlU6iMiaOmUntibsCTZtgFl/D1
HpI+bfQ5ubwHc0ygxTCKGPqQKOl0cXxpzsvAIr0z9k9MD6WHl0s2m7QwGehEW689
qHMQs4y1xe4sT+igg29/6c7XYGTtefm5ojDMC/cSjjf7FiR01n0JltIHPsxRhkTs
iHm3rfYJV37K5RQk9lXeQT7lqY1RQrn2JhzX/3cXFatHzws4J+4CEbEH8/iAryg8
NO5qDSAOrVFqYh06tFlUerGXIN9d4M+oVmFg1Bmrf5/p4iLcTi2gsO6Q/36Vbu9H
AWx/LR5jJlVc5OedkmeNxeETI/f0vf+TUQgHaJ/D8M/Iof0Eu6BMzaxEclkdvnZf
3Yatzbvrope30TWLnhr19zQcc/fkW1AjkKfbsA62pNDIQKNwd5Xitvzmv0bhbf88
vyGyZv5MlwEJsGDo6opdA7e21Tj9tN7Lo5mSiqyAcozH8GuUQrCn8lAvRF+IfqIW
v/Vr4r2XfdeCLRDjA1S+bzujeLLmLvI1Mt/SFNshx8ZsDNO0D2IJNHF6vT1fB278
NNWmn+F0U5eKG9NIRa4xW1B58PvGyWv6WKFYiunWheTqJelePVO2oZVs/htAgIuO
K6ccvUOGbu8HYLt7AfrxAk4LllUgt4kryZmKqddoj+SfuwtiWHj6pTveEm2fna6n
8ggU6Em0KmdEESGKdBPzSZ7FMYx0XUszHAG340ReaYxtriS6yRohdboMLDMSums9
WM2cER93ev4xgNKCIMpJvdET5l6mkbs/1zwhwl15NS9xW7/EUxokUp+LPKMNMCqn
2ZjKBR3fEuL7565WhjCOxboO5wGQgF9rNqikkz1EEuwNanPnOL24ZxggXmbOufm2
O/mVeNQUrxBvKBcApycqwCuAPOjZhQ59tz3ajrZcWj7yv2OaI1yrxMQuhv4o9fHl
WZ+sicf8IL8xYPJOoFpseG2dqVHiJTrcie388kAPwnND8NF2wMc/0erxVlf1cNoj
YnThjtJ5tjTus0TPrX1zUmrDT/W1ZxBpPv9C/wcTgg4Q1tKNxmzExgPQybharc0q
wQ7tBBv5yTuTZ1LfIp1XU32BAOLCD0kZOgXNa9es4EDTG6A+AkYCLaGt6zBiQc5d
La6F1dr7IsAt4Sn7LAiiMhNVJdESwNJZQLQMnCBr2osPz+HCsGCB68UncF55qQCa
sXsUnov6fVzHqhHMUUFOSSq1mBmqhnnJG39wIH+Ud24ZhTDV2/+GL/rOPehpxg81
GoQI/Ugc/l/LSb5iRGRrj8Pfq/a2bgeqa0FevUCuKcfvD3aRSlmknqTI6zvBcf28
BbXoXM8jSSErATgDgTMPXZRJCPEUjpv3FLVQmniMKH/B0JhKvmqPpw77FuUDPPaM
N8v7x7XyRaMNvmvgouVlobc+jyiohxrZYber7ieBgRul4wACGzD02ULimxg1qCYY
lQIPPw3X7FDR1yn6KDeVnl4dsR12a+8ieZ/Exr7DgqZRk56CdZ0kHRhLeX9WMDxP
E7p/NSWzp0eG0znLN7+XvMUYdlFe6rJRBk+l3WsXdlr6hkntLfXcIiH1bveTiSIu
1pcpapJxMmf2IGR3b/BDUZBMtEU+b1cZ3vjTysGC8edqe4ZERtVrPuqx3X7dJA5a
PkHnnb6G1+gyLVX9HE2YESA7qNvdr4KsSts8wU7Clmam1FMxKzq3jBP9fxKrKqP8
ApE4M/uYhl7pB4fJGJMKntLRLFKrKfkPg34Gg1ESX0MIgUliE7iA0VE3AE8W2Gca
A/UTIsucQ4UhxQgmJsUVHno3R+/5xiSEbT8pNS1rcVQFV3T0olYo9wXCWkDeZF9R
e/QsLLLRkzNj2hkZhS1dqFaOYSqldLa5XP2jHnjT37K3s+pP5DvWczvYm/9wLv25
oKq2xzVzvPGMB/MynMlthKGwwvD8Jav1YkvBl3by9L9CWJpdk3S+ZrBGJ7LyhLFf
TlPNJRv+z5cx/3G/xR7EVt96UXV5NFFqjgTNbFOdAYDC3R+IZuopr4iwvTbjDsTf
6iOBAZEDDrRozMXrubcmkGZF+BoCbs3ci+80lJZ3rMiLJU4BIDC6FshqTFsK63RH
nNbbdyPFYDY3VXKMCZDAZEcYVUM8MDSBmKZF7UfqA8xo/SzGub4PSoa4N6FdldWG
7t6oC3xgtbkMCtyBoSwGge8yoSPSkNI0aBH5APmtNuu3/Tyd3h0zFcfqf2jU82Gj
AsWVEe7skj41SvWJA0srfWX18gSJRekhgwNuKkUw3NUH/2uah8VW5shAZQs/w7OS
dVy3ra8iEcv8hWgNOlMym9GkYD/VNx+F83LYnPOXyLX48HrUmEYwHlSR8vDRQJA7
sOR5aKBxpk6S4vbnaEJpqwVLP/bJPLcXuLZm4imW5Lqutx26LK7ACN7OJDHQ7rMQ
RlQK/oKRoZy9tMsvwT14JMJKzoDwxMJhnDXU/CQOFo4xZCohddq8RCDNZ/2ICuXs
YfbjG6ajqZlzJHM0Jwc4cxcDOJvbSydHMM259KYWmscLWnMAER83k6Q24cro4BUy
/nUGTYuBgq1LRpd+3MwgJcLyGBNdcVOS4USh4QpSj14NK85ALVu1HG2HiozNnxEp
/e0MTbnwld+lWL3pvO1A/y65kjAikHMY8wQCf7chrRijt0iSIpgwgQpl1kWCu5tu
CaBi7AAg5gTd8tcnsPsEUjbMgoMn0/VKtQc/MCvvyJ42MVPAjZITnrYcyScUewtQ
yr2/lynzqxk/IQCaDaHdvoHD0PocomHZI9TbzUfzpBHA6ZXnmRrISHgbTAR8JEBJ
pHjj79ofbm/ZW+eaqOKHoUkPmCEmwh02d17Q6hmf7Q5CdgkL8uDrfnnuRx1s8z+b
WTlDxHs15knOFkRMjmAS7nQGdmpEQ6BeV97h0VV0bggaAi6xSGrRJT/y+4Pj/zTq
EWi4+Y2SsuzeOfIxVU4bF5ToKalMzG21ds5wHNb82Xqlz5PIFI4DBYlIA/bq3s+m
2DN3Zxj55wFIqf5Ih/A0cdWcsfXzN0SvNn5CbcJ4LBIPX/L999boVIYSbjOP1jb2
cidsfsWThVo/c5JYgMpPpiUD22c5MzW3wPXdANsunNeRATyjYPAMKN3dMdhhX+Gh
7MLrgYwwMLdJK6MqZsBO9hENxVLR0fOINsZUu0rNpKPkWt/J350Itmi4uEx2DIc+
FThB+GO7hpddsF3mJ5GQgBTVpQwquyQepC6rujQSpQTmfz3FADD/SE+fV8xhK/UP
eKrsVjgnGDISdKgGg/WzsiPvQh8lNPansiA6cxxZEooDk3gx3wjmE3evvMAv8o5U
3OVNBGymJo9W3POVzNiZkLlgzhA6uZMPACG26Vd6vqfyZds9tEXYGHRs8GhC75w2
uSgxMjww0dbGwEQ+D0xDXmaT3WP+c0YMkTQKaRUSumNbCpFevVDYIuKXrVxCYu/C
cBfKcGWyYtWk52LXxyJ5zI9nMnfTmgLa1O+N939UXDXztZ6Gw3Xe3KlCNtqSMcgK
uI95B1IZCZNzaGvS2sGfo8QRgYJHu6pVVXHsaBB3QrEkfkdGwz7sR4QI+RT4/tTM
IMIe1QqMwD/74PCKhC/65EYgIvaFLLJZNPELpKqWoLWqfeIyGmVrf+gkxocKii1H
JH91Gc5rnB7OQT6yXWAS6fQSaptVb7cp6TDmuAdpirbDNpTxs2r/D6zeapl3lxAD
/psrm+Lz908ZqElMs+R1idSQofeK+bb1uVqZhvnaPzCPvspvKwnA5cEKF4TWwErW
iZ1c79a0Kpw0ZX6Mr7azJIJKa0PopF7/6n8g2rI8VP6eP3QyF5cI2wYrmtXsAsQX
mcpw/qB2P46EJsZOiuDDcIYD36ErIl/y5DQTlOiv33xoYpnhw7W1Y7axTqdjyl0p
aeflqK4Wv2VRABFqIcjafgopg1m/FC7z0mriGLuC1HQFHzFU1dHPFvco0Gf2+aIT
qdz6Ty8C0xaNRqYkU7H7vnsXN+yyUqcI5+59cEqrlXduMqO/76xUdgUZd8b7e9HT
PeOk3rBO0a2juF3G2Ct4bBOovFY5gAG0VG83U1IwqPWwt3TpicP5uDQuybKhwPGf
DuUXbBxpp0Bpxmh5oWJfVYF/TPWN60gADXuNfRtKcCDjgevkJ9vex3mpONd6udQv
LlxyUb6L7gCZFuv37mWyYS8+yIgJza+CU8oIWXIQMDXne/vQWDsYEIPysNN/njiZ
LTG9xlIDYe2lTiPv0leAmlVoY1WeE4eVM44ICgOD/rhauP25fAK4mu9KCmG6bU2y
08G+FTOHxpnhV0dh/Xyz9LI1z/VBUL/x1UhNK5bOybJO+pwBwNiK9NCq+TgARRcL
Ag+uybLmiZIUbda2jey8+L5mlV7Y5zM4wRrchRZhTb9Z2Ef3XJMCsSNC0hwvwui6
gbyok7jPJV3ehF2mlBYwZFbMvXKJkhsylS/EJRBuDXemDKGnajkjXrjrh/opZ1YB
Q1S1TfDg2V7CmKYh/YRvH5n3w3nO6vJeXUo7Scj4+KkeTKd8uPW99h6n2zaWJ/KZ
hQB4YXpdkCHTfiCVXUYW8uypARsdiajCLQmIfvK3fk+VGfOBH+tToGqFYaXtHsMp
MkfPndnA/k1vXnQDlubkS3+zKpJP2H+BytplOPl7ZhSOdmFy3MWSpHL9gERkGx8n
EpTG+6sXUnpSYDR8N3TMvXbus97jlGtod66JxbIgwtvrChDB1fmpB7SJG/ahBO6Y
VlEH9uR9bxU7hX/1D6U63CwOTu4CiOJhb2mOYjjuxMM4O5DZsjsl5aeZopFoilV/
siUzJQS8ruEZx+b4IjCBXqj5xHur3uqjU9u6hdlqVS1DxgK2Dt+Nb9Cx0e33p3aC
zrYdcGa9r8a1itcnHRAFD7X/QcQuqvOT3zSSofLnQJsF0/gLSKRZltfeeGFv7SH6
T1uge2yABl7MfJguRFfPd7+ASuu+4H8CX7SaX4eihUpNxsy1hgLAw/upnBgbgHd7
J2XmvkOzXQlZyj5yyzFEh6mCX/Wplra9r/o/aT8xQA2xEyPcCQLWrbmUMx7d/HAS
X1/bLxJmR8Omn700xHe3QZTCgSQ/b7PjExsJ6RyRVJJ7PqSu0Vkx4EAFiaSxQU8I
MPbgbJFAETcV4ZYsGIzjpSl7xoR39V+nUhCVNSAVhEn7Caf1ZyHJzQynZxA48sWT
/i1OFs70wB4X5UfUD3u6e2W5OLFDbAnKkPuGTasgCoS2gjU9WYl5zMfSeNBp/O1k
WXRIi7FzzJfJ3v/o7hhpl2nsbAzHTzT5vf/GAI2T04nSde7U6FA2CrJqymMuw8sS
e2HxpyXrh84m0Jh03smugIYWDDLwSNg/djen0uNHVGjpnHvGXyExChHHmY6uDIE/
3ZUR9DdHVBxwudJrpZckKJ9uiPSPzgccbFQYRiMMdRugFQ/LoFaXJOMNQKzooz2t
DRzTyNpLvp9FJBH9bj9+abzgTA7GBO+6AqBAqk4ZN134bDtMfI9P3O/TBYrTOJYi
SA+ggtVYH+CNlMONN71sw2FdgYHUIZQUqDbys86n+UXp7PRiZz9WZza7k709RpDx
brQXY4EZjY/DRXfo4RQd+7E1A6vr1W1eZsS9zUmP6KZh8N+y8SZYzMROSE0Eqzx+
+mNidIBraGjcmqToBL87ufAb4ii+/WZMzwp8CuFSHxEGUxDPZpzHYTluIQIDP40d
ydwvJshXXGqk2nBnc5mUSab4W8iAsiSkjvps2jWT3x4mOE4Nsd/wq9feC6sxitup
0nEVnqLKN/PF3E98b33q1TeBDr7URyeBdmbLcEewytuRJxq2yg1w4w6yAVC6vZrb
RZCHusemZb8Wdb5K4e993goB1KtYF2dCyS+HTVibrEJVaWGGdgzLchri+jT/wSDp
oudTeJOA4XneNoJnZgL0sIdDx0tjTNdFEpok9f6h3tDMPxFAs8D13P53GzYluJg8
TtJNLTA5Uyvc4zIT/6k1OlX2jibUOAF0/h3OqQVvIwAcJASpRQr50eug5rGg0QaA
sMeqhgOXcoH84/Auoyl9cvX7hOMXFSETfxgUabIeZv10s1bZSfdWI5e/7EjyYIHV
tRV8swuee1MWESNQaPuqZ6178yWtQdgd6yQQ9tbPBCOQfIT+rpUFokc4JOhuzrX0
x1zWwgFiH3K+CMbskBrzTUA6Fz0AeSKhDMNX/Ku2Vi12ez56UMhwgohlfohxyt3L
kSXzsdlyCYszBzaNEdBnpYOoXZErj5eWnahFtaE/Y9VtmZf2fl9dxuk/m8L2Vk9t
bbLIpJ0G4nMrmQrsOozV1LQJtxIHRlQYbl2KNCB6u9T68Lb3c7mE07GlpPUJImAX
gG39gC/ddyoRBfATELnsYAkMHXkAcFEunzyRZQiqoKBFPWfgmP/g0JHQHzGGm/Hu
kgeD32z+TlLDQjLf75NIQt9Keno2w/jp+2+8sbrXDXVwnqjpxiS57CB9dve4FWJG
ssFEAXcTdVQvSn45auI+Vz6WZPwNwtgI3i61sF8C3zg+UtWIh+6pJHjGHLw1vvpl
pQ9FydR537cX6BDa0LJAgJ4+3yUKKEvfMtVC4jltgNhpWcG1D2tMozSN1gdu/lKI
2ji08GlmgsneCJgGWOuHM2wmUm9sAm8cfPygOqXbiDYLXyn2B53FcsZgWXBX/uyc
Z6GwyApZv1OlwdtUG3oyf32swZpTVAbPw6IIds1ICEmqsDQDZ/IOwnsv1/TiyUoS
vtaBPo9De3yp6R8ELQhPjNnngTMxh+OVu7qhB+XaiFs=
//pragma protect end_data_block
//pragma protect digest_block
IaCqQvdrcyahbwCySguXdNHAtb4=
//pragma protect end_digest_block
//pragma protect end_protected
