
`define CYCLE_TIME 20.0
`define SEED_NUMBER 38524879
`define PATTERN_NUMBER 100
`define DEBUG_MODE 1 // This will generate a "process.txt" file for debugging

module PATTERN(
  // Output signals
  output reg clk, rst_n, in_valid, in_valid2,
  output reg [7:0] image, template,
  output reg [1:0] image_size,
  output reg [2:0] action,
  // Input signals
	input out_valid, out_value
);
// ========================================
// clock
// ========================================
real CYCLE = `CYCLE_TIME;
always	#(CYCLE/2.0) clk = ~clk;
// ========================================
// integer & parameter
// ========================================
integer SEED;
integer pat_count, act_count;
integer f_img, f_img_h;
integer i, j, k, l, m;
integer exe_latency, total_latency;
// ========================================
// wire & reg
// ========================================
reg [7:0] test_R[0:15][0:15], test_G[0:15][0:15], test_B[0:15][0:15];
reg [7:0] gray_M[0:15][0:15], gray_A[0:15][0:15], gray_W[0:15][0:15];
reg [7:0] test_template[0:2][0:2];
reg [1:0] test_size;
integer img_size;
reg [3:0] test_action[0:7];
integer action_num;
reg [7:0] temp[0:15][0:15], temp1[0:15][0:15];
integer golden_size;
reg [19:0] golden_out[0:15][0:15];
reg [19:0] rec_out[0:15][0:15];

reg [7:0] a0, a1, a2, a3, a4, a5, a6, a7, a8;
reg check;
//================================================================
// design
//================================================================
initial begin
  reset_task;
  for(pat_count = 0; pat_count < `PATTERN_NUMBER; pat_count = pat_count + 1) begin
    input_img_task;
    for(act_count = 0; act_count < 8; act_count = act_count + 1) begin
      input_action_task;
      ans_gen_task;
      wait_task;
      check_task;
    end
  end
  YOU_PASS_task;
end

always @(negedge clk) begin
  if(out_valid === 1'b0 && out_value !== 1'b0) begin : OUT_RESET_CHECK
    fail_task;
    $display("--------------------------------------------------");
    $display("                      FAIL!!                      ");
    $display("      Output must be 0 when out_valid is low      ");
    $display("--------------------------------------------------");
    repeat(5) @(negedge clk);
    $finish;
  end
  if(in_valid === 1'b1 && out_valid === 1'b1) begin : OVERLAP_CHECK
    fail_task;
    $display("--------------------------------------------------");
    $display("                      FAIL!!                      ");
    $display("   in_valid and out_valid cannot be high at once  ");
    $display("--------------------------------------------------");
    repeat(5) @(negedge clk);
    $finish;
  end
end
//---------------------------------------------------------------------
//   Task
//---------------------------------------------------------------------
task reset_task;
  SEED = `SEED_NUMBER;
  rst_n = 1'b1;
  in_valid = 1'b0;
  in_valid2 = 1'b0;
  image = 8'dx; template = 8'dx; image_size = 2'dx; action = 3'dx;

  total_latency = 0;

  force clk = 'b0;
  #(CYCLE * ($random(SEED) % 'd3 + 'd1)); rst_n = 'b0;
  #(CYCLE * 0.75);

  if(out_valid !== 1'b0 || out_value !== 1'b0) begin : RESET_CHECK
    fail_task;
    $display("--------------------------------------------------");
    $display("                      FAIL!!                      ");
    $display("           Output must be 0 after reset           ");
    $display("--------------------------------------------------");
      #(CYCLE * 5);
    $finish;
  end

  #(CYCLE * 0.25); rst_n = 'b1;
  #(CYCLE); release clk;
  repeat(3) @(negedge clk);
endtask

task input_img_task;
  repeat($random(SEED) % 'd3 + 'd1) @(negedge clk);
  if(pat_count == 0)
    test_size = 2'd0;
  else if(pat_count == 1)
    test_size = 2'd1;
  else if(pat_count == 2)
    test_size = 2'd2;
  else
    test_size = $random(SEED) % 'd3;
  case(test_size)
    2'd0: img_size = 4;
    2'd1: img_size = 8;
    2'd2: img_size = 16;
  endcase
  for(i = 0; i < 9; i = i + 1)
    test_template[i / 3][i % 3] = $random(SEED) % 'd256;

  in_valid = 1'b1;
  k = 0;
  for(i = 0; i < img_size; i = i + 1) begin
    for(j = 0; j < img_size; j = j + 1) begin
      image_size = (i == 0 && j == 0) ? test_size : 2'dx;
      test_R[i][j] = $random(SEED) % 'd256;
      test_G[i][j] = $random(SEED) % 'd256;
      test_B[i][j] = $random(SEED) % 'd256;

      image = test_R[i][j];
      template = (k < 9) ? test_template[k / 3][k % 3] : 8'dx;
      k = k + 1;
        @(negedge clk);
      image_size = 2'dx;
      image = test_G[i][j];
      template = (k < 9) ? test_template[k / 3][k % 3] : 8'dx;
      k = k + 1;
        @(negedge clk);
      image = test_B[i][j];
      template = (k < 9) ? test_template[k / 3][k % 3] : 8'dx;
      k = k + 1;
        @(negedge clk);
    end
  end
  in_valid = 1'b0;
  image = 8'dx; template = 8'dx; image_size = 2'dx;
    @(negedge clk);
endtask

task input_action_task;
  repeat($random(SEED) % 'd3 + 'd1) @(negedge clk);
  action_num = $random(SEED) % 'd7 + 'd2;
  test_action[0] = $random(SEED) % 'd3;
  for(i = 1; i < action_num - 1; i = i + 1)
    test_action[i] = $random(SEED) % 'd4 + 'd3;
  test_action[action_num - 1] = 3'd7;

  in_valid2 = 1'b1;
  i = 0;
  repeat(action_num) begin
    action = test_action[i];
    i = i + 1;
      @(negedge clk);
  end
  in_valid2 = 1'b0;
  action = 3'dx;
    @(negedge clk);
  exe_latency = 1;
endtask

task ans_gen_task;
  if(`DEBUG_MODE) begin
    f_img = $fopen("process.txt", "w");
    f_img_h = $fopen("process_hex.txt", "w");
    $fdisplay(f_img, " Image(R)");
    $fdisplay(f_img_h, " Image(R)");
    print_array(f_img, img_size, test_R);
    print_hex(f_img_h, img_size, test_R);
    $fdisplay(f_img, " Image(G)");
    $fdisplay(f_img_h, " Image(G)");
    print_array(f_img, img_size, test_G);
    print_hex(f_img_h, img_size, test_G);
    $fdisplay(f_img, " Image(B)");
    $fdisplay(f_img_h, " Image(B)");
    print_array(f_img, img_size, test_B);
    print_hex(f_img_h, img_size, test_B);
    $fdisplay(f_img, "Template");
    $fwrite(f_img, "  ");
    for(i = 0; i < 3; i = i + 1) $fwrite(f_img, " %3d", i);
    $fwrite(f_img, "\n----");
    for(i = 0; i < 3; i = i + 1) $fwrite(f_img, "----");
    $fwrite(f_img, "\n");
    for(i = 0; i < 3; i = i + 1) begin
      $fwrite(f_img, "%2d| ", i);
      for(j = 0; j < 3; j = j + 1) begin
        $fwrite(f_img, "%3d ", test_template[i][j]);
      end
      $fwrite(f_img, "\n");
    end
    $fdisplay(f_img_h, "Template");
    $fwrite(f_img_h, "  ");
    for(i = 0; i < 3; i = i + 1) $fwrite(f_img_h, " %2d", i);
    $fwrite(f_img_h, "\n----");
    for(i = 0; i < 3; i = i + 1) $fwrite(f_img_h, "---");
    $fwrite(f_img_h, "\n");
    for(i = 0; i < 3; i = i + 1) begin
      $fwrite(f_img_h, "%2d| ", i);
      for(j = 0; j < 3; j = j + 1) begin
        $fwrite(f_img_h, "%2h ", test_template[i][j]);
      end
      $fwrite(f_img_h, "\n");
    end
    for(j = 0; j < img_size; j = j + 1) begin
      for(k = 0; k < img_size; k = k + 1) begin
        gray_M[j][k] = (test_R[j][k] > test_G[j][k]) ? test_R[j][k] : test_G[j][k];
        gray_M[j][k] = (gray_M[j][k] > test_B[j][k]) ? gray_M[j][k] : test_B[j][k];
      end
    end
    $fdisplay(f_img, "\nGrayscale - Max");
    $fdisplay(f_img_h, "\nGrayscale - Max");
    print_array(f_img, img_size, gray_M);
    print_hex(f_img_h, img_size, gray_M);
    for(j = 0; j < img_size; j = j + 1) begin
      for(k = 0; k < img_size; k = k + 1) begin
        gray_A[j][k] = (test_R[j][k] + test_G[j][k] + test_B[j][k]) / 3;
      end
    end
    $fdisplay(f_img, "Grayscale - Average");
    $fdisplay(f_img_h, "Grayscale - Average");
    print_array(f_img, img_size, gray_A);
    print_hex(f_img_h, img_size, gray_A);
    for(j = 0; j < img_size; j = j + 1)
      for(k = 0; k < img_size; k = k + 1)
        gray_W[j][k] = (test_R[j][k] >> 2) + (test_G[j][k] >> 1) + (test_B[j][k] >> 2);
    $fdisplay(f_img, "Grayscale - Weighted");
    $fdisplay(f_img_h, "Grayscale - Weighted");
    print_array(f_img, img_size, gray_W);
    print_hex(f_img_h, img_size, gray_W);
    $fwrite(f_img, "\nAction :");
    $fwrite(f_img_h, "\nAction :");
    for(i = 0; i < action_num - 1; i = i + 1) begin
      $fwrite(f_img, "%2d ->", test_action[i]);
      $fwrite(f_img_h, "%2d ->", test_action[i]);
    end
    $fdisplay(f_img, "%2d\n", test_action[action_num - 1]);
    $fdisplay(f_img_h, "%2d\n", test_action[action_num - 1]);
  end
  golden_size = img_size;
  for(i = 0; i < action_num; i = i + 1) begin
    case(test_action[i])
      // Grayscale - Max
      3'd0: begin
        for(j = 0; j < golden_size; j = j + 1) begin
          for(k = 0; k < golden_size; k = k + 1) begin
            temp[j][k] = (test_R[j][k] > test_G[j][k]) ? test_R[j][k] : test_G[j][k];
            temp[j][k] = (temp[j][k] > test_B[j][k]) ? temp[j][k] : test_B[j][k];
          end
        end
        if(`DEBUG_MODE) $fdisplay(f_img, "Action 0 (Grayscale - Max)");
        if(`DEBUG_MODE) $fdisplay(f_img_h, "Action 0 (Grayscale - Max)");
        if(`DEBUG_MODE) print_array(f_img, golden_size, temp);
        if(`DEBUG_MODE) print_hex(f_img_h, golden_size, temp);
      end
      // Grayscale - Average
      3'd1: begin
        for(j = 0; j < golden_size; j = j + 1) begin
          for(k = 0; k < golden_size; k = k + 1) begin
            temp[j][k] = (test_R[j][k] + test_G[j][k] + test_B[j][k]) / 3;
          end
        end
        if(`DEBUG_MODE) $fdisplay(f_img, "Action 1 (Grayscale - Average)");
        if(`DEBUG_MODE) $fdisplay(f_img_h, "Action 1 (Grayscale - Average)");
        if(`DEBUG_MODE) print_array(f_img, golden_size, temp);
        if(`DEBUG_MODE) print_hex(f_img_h, golden_size, temp);
      end
      // Grayscale - Weighted
      3'd2: begin
        for(j = 0; j < golden_size; j = j + 1)
          for(k = 0; k < golden_size; k = k + 1)
            temp[j][k] = (test_R[j][k] >> 2) + (test_G[j][k] >> 1) + (test_B[j][k] >> 2);
        if(`DEBUG_MODE) $fdisplay(f_img, "Action 2 (Grayscale - Weighted)");
        if(`DEBUG_MODE) $fdisplay(f_img_h, "Action 2 (Grayscale - Weighted)");
        if(`DEBUG_MODE) print_array(f_img, golden_size, temp);
        if(`DEBUG_MODE) print_hex(f_img_h, golden_size, temp);
      end
      // Max pooling
      3'd3: begin
        if(golden_size == 4) begin
          for(j = 0; j < 4; j = j + 1)
            for(k = 0; k < 4; k = k + 1)
              temp[j][k] = temp1[j][k];
        end else begin
          for(j = 0; j < golden_size; j = j + 2) begin
            for(k = 0; k < golden_size; k = k + 2) begin
              temp[j / 2][k / 2] = (temp1[j][k] > temp1[j + 1][k]) ? temp1[j][k] : temp1[j + 1][k];
              temp[j / 2][k / 2] = (temp[j / 2][k / 2] > temp1[j][k + 1]) ? temp[j / 2][k / 2] : temp1[j][k + 1];
              temp[j / 2][k / 2] = (temp[j / 2][k / 2] > temp1[j + 1][k + 1]) ? temp[j / 2][k / 2] : temp1[j + 1][k + 1];
            end
          end
          golden_size = golden_size / 2;
        end
        if(`DEBUG_MODE) $fdisplay(f_img, "Action 3 (Max pooling)");
        if(`DEBUG_MODE) $fdisplay(f_img_h, "Action 3 (Max pooling)");
        if(`DEBUG_MODE) print_array(f_img, golden_size, temp);
        if(`DEBUG_MODE) print_hex(f_img_h, golden_size, temp);
      end
      // Negative
      3'd4: begin
        for(j = 0; j < golden_size; j = j + 1)
          for(k = 0; k < golden_size; k = k + 1)
            temp[j][k] = 'd255 - temp1[j][k];
        if(`DEBUG_MODE) $fdisplay(f_img, "Action 4 (Negative)");
        if(`DEBUG_MODE) $fdisplay(f_img_h, "Action 4 (Negative)");
        if(`DEBUG_MODE) print_array(f_img, golden_size, temp);
        if(`DEBUG_MODE) print_hex(f_img_h, golden_size, temp);
      end
      // Horizontal Flip
      3'd5: begin
        for(j = 0; j < golden_size; j = j + 1)
          for(k = 0; k < golden_size; k = k + 1)
            temp[j][k] = temp1[j][golden_size - k - 1];
        if(`DEBUG_MODE) $fdisplay(f_img, "Action 5 (Horizontal Flip)");
        if(`DEBUG_MODE) $fdisplay(f_img_h, "Action 5 (Horizontal Flip)");
        if(`DEBUG_MODE) print_array(f_img, golden_size, temp);
        if(`DEBUG_MODE) print_hex(f_img_h, golden_size, temp);
      end
      // Image Filter
      3'd6: begin
        for(j = 0; j < golden_size; j = j + 1) begin
          for(k = 0; k < golden_size; k = k + 1) begin
            a0 = (j == 0 && k == 0) ? temp1[j][k] : 
                 (j == 0) ? temp1[j][k - 1] : 
                 (k == 0) ? temp1[j - 1][k] : temp1[j - 1][k - 1];
            a1 = (j == 0) ? temp1[j][k] : temp1[j - 1][k];
            a2 = (j == 0 && k == golden_size - 1) ? temp1[j][k] : 
                 (j == 0) ? temp1[j][k + 1] : 
                 (k == golden_size - 1) ? temp1[j - 1][k] : temp1[j - 1][k + 1];
            a3 = (k == 0) ? temp1[j][k] : temp1[j][k - 1];
            a4 = temp1[j][k];
            a5 = (k == golden_size - 1) ? temp1[j][k] : temp1[j][k + 1];
            a6 = (j == golden_size - 1 && k == 0) ? temp1[j][k] : 
                 (j == golden_size - 1) ? temp1[j][k - 1] : 
                 (k == 0) ? temp1[j + 1][k] : temp1[j + 1][k - 1];
            a7 = (j == golden_size - 1) ? temp1[j][k] : temp1[j + 1][k];
            a8 = (j == golden_size - 1 && k == golden_size - 1) ? temp1[j][k] : 
                 (j == golden_size - 1) ? temp1[j][k + 1] : 
                 (k == golden_size - 1) ? temp1[j + 1][k] : temp1[j + 1][k + 1];
            temp[j][k] = median(a0, a1, a2, a3, a4, a5, a6, a7, a8);
          end
        end
        if(`DEBUG_MODE) $fdisplay(f_img, "Action 6 (Image Filter)");
        if(`DEBUG_MODE) $fdisplay(f_img_h, "Action 6 (Image Filter)");
        if(`DEBUG_MODE) print_array(f_img, golden_size, temp);
        if(`DEBUG_MODE) print_hex(f_img_h, golden_size, temp);
      end
      // Cross Correlation
      3'd7: begin
        for(j = 0; j < golden_size; j = j + 1) begin
          for(k = 0; k < golden_size; k = k + 1) begin
            golden_out[j][k] = 0;
            for(l = -1; l < 2; l = l + 1) begin
              for(m = -1; m < 2; m = m + 1) begin
                if(j + l >= 0 && j + l < golden_size && k + m >= 0 && k + m < golden_size)
                  golden_out[j][k] = golden_out[j][k] + temp1[j + l][k + m] * test_template[l + 1][m + 1];
              end
            end
          end
        end
        if(`DEBUG_MODE) begin
          $fwrite(f_img, "Action 7 (Cross Correlation)\n   ");
          for(j = 0; j < golden_size; j = j + 1) $fwrite(f_img, " %7d", j);
          $fwrite(f_img, "\n----");
          for(j = 0; j < golden_size; j = j + 1) $fwrite(f_img, "--------");
          $fwrite(f_img, "\n");
          for(j = 0; j < golden_size; j = j + 1) begin
            $fwrite(f_img, "%2d| ", j);
            for(k = 0; k < golden_size; k = k + 1) begin
              $fwrite(f_img, "%7d ", golden_out[j][k]);
            end
            $fwrite(f_img, "\n");
          end
          $fwrite(f_img, "\n");
          $fwrite(f_img_h, "Action 7 (Cross Correlation)\n   ");
          for(j = 0; j < golden_size; j = j + 1) $fwrite(f_img_h, " %5d", j);
          $fwrite(f_img_h, "\n----");
          for(j = 0; j < golden_size; j = j + 1) $fwrite(f_img_h, "------");
          $fwrite(f_img_h, "\n");
          for(j = 0; j < golden_size; j = j + 1) begin
            $fwrite(f_img_h, "%2d| ", j);
            for(k = 0; k < golden_size; k = k + 1) begin
              $fwrite(f_img_h, "%5h ", golden_out[j][k]);
            end
            $fwrite(f_img_h, "\n");
          end
          $fwrite(f_img_h, "\n");
        end
      end
    endcase
    for(j = 0; j < golden_size; j = j + 1)
      for(k = 0; k < golden_size; k = k + 1)
        temp1[j][k] = temp[j][k];
  end
  if(`DEBUG_MODE) $fclose(f_img);
  if(`DEBUG_MODE) $fclose(f_img_h);
endtask

function reg [7:0] median;
  input reg [7:0] a0, a1, a2, a3, a4, a5, a6, a7, a8;
  reg [7:0] sorted[0:8];
  begin
    sorted[0] = a0; sorted[1] = a1; sorted[2] = a2;
    sorted[3] = a3; sorted[4] = a4; sorted[5] = a5;
    sorted[6] = a6; sorted[7] = a7; sorted[8] = a8;
    sorted.sort();
    median = sorted[4];
  end
endfunction

task print_array;
  input integer file, size;
  input reg [7:0] array[0:15][0:15];
  integer p, q;
  begin
    $fwrite(file, "    ");
    for(p = 0; p < size; p = p + 1) $fwrite(file, "%3d ", p);
    $fwrite(file, "\n----");
    for(p = 0; p < size; p = p + 1) $fwrite(file, "----");
    $fwrite(file, "\n");
    for(p = 0; p < size; p = p + 1) begin
      $fwrite(file, "%2d| ", p);
      for(q = 0; q < size; q = q + 1) begin
        $fwrite(file, "%3d ", array[p][q]);
      end
      $fwrite(file, "\n");
    end
    $fwrite(file, "\n");
  end
endtask

task print_hex;
  input integer file, size;
  input reg [7:0] array[0:15][0:15];
  integer p, q;
  begin
    $fwrite(file, "    ");
    for(p = 0; p < size; p = p + 1) $fwrite(file, "%2d ", p);
    $fwrite(file, "\n----");
    for(p = 0; p < size; p = p + 1) $fwrite(file, "---");
    $fwrite(file, "\n");
    for(p = 0; p < size; p = p + 1) begin
      $fwrite(file, "%2d| ", p);
      for(q = 0; q < size; q = q + 1) begin
        $fwrite(file, "%2h ", array[p][q]);
      end
      $fwrite(file, "\n");
    end
    $fwrite(file, "\n");
  end
endtask

task wait_task;
  while(out_valid !== 1'b1) begin
    exe_latency = exe_latency + 1;
    if(exe_latency == 5000) begin : TIMEOUT_CHECK
      fail_task;
      $display("--------------------------------------------------");
      $display("                      FAIL!!                      ");
      $display("       Execution timeout (over 5000 cycles)       ");
      $display("--------------------------------------------------");
      repeat(5) @(negedge clk);
      $finish;
    end
      @(negedge clk);
  end
endtask

task check_task;
  i = 0; j = 0; check = 0;
  repeat(golden_size ** 2) begin
    for(k = 19; k >= 0; k = k - 1) begin
      rec_out[i][j][k] = out_value;
      if(out_valid !== 1'b1) begin
        fail_task;
        $display("--------------------------------------------------");
        $display("                      FAIL!!                      ");
        $display("        out_valid should high consecutively       ");
        $display("--------------------------------------------------");
        repeat(5) @(negedge clk);
        $finish;
      end
        @(negedge clk);
    end
    if(rec_out[i][j] !== golden_out[i][j]) begin
      check = 1;
    end
    j = (j == golden_size - 1) ? 0 : j + 1;
    i = (j == 0) ? i + 1 : i;
  end
  if(out_valid !== 1'b0) begin
    fail_task;
    $display("--------------------------------------------------");
    $display("                      FAIL!!                      ");
    $display("        out_valid must be low after output        ");
    $display("--------------------------------------------------");
    repeat(5) @(negedge clk);
    $finish;
  end
  if(check) begin
    fail_task;
    $display("--------------------------------------------------");
    $display("                      FAIL!!                      ");
    $display("         Output does not match with golden        ");
    $display("==================================================");
    $display("  Golden:");
    for(i = 0; i < golden_size; i = i + 1) begin
      for(j = 0; j < golden_size; j = j + 1) begin
        $write(" %7d", golden_out[i][j]);
      end
      $display("");
    end
    $display("  Yours:");
    for(i = 0; i < golden_size; i = i + 1) begin
      for(j = 0; j < golden_size; j = j + 1) begin
        if(rec_out[i][j] !== golden_out[i][j])
          $write("\033[38;5;196m %7d\033[0m", rec_out[i][j]);
        else
          $write(" %7d", rec_out[i][j]);
      end
      $display("");
    end
    $display("\n--------------------------------------------------");
    repeat(5) @(negedge clk);
    $finish;
  end
  $display("\033[38;5;123mPATTERN NO.%4d\033[0;38;5;150m ACTION NO.%2d PASS!!\033[0;32m EXECUTION CYCLE :%4d\033[m", pat_count, act_count, exe_latency);
  total_latency = total_latency + exe_latency;
endtask

task YOU_PASS_task;
  $display("\033[0m                                                \033[38;2;255;255;255m$\033[38;2;250;252;252m@\033[38;2;255;255;255m$$\033[0m                                                                             \033[0m");
  $display("\033[0m                                                \033[38;2;255;255;255m$\033[38;2;255;249;234mB\033[38;2;224;215;202m*\033[38;2;247;248;251m@\033[38;2;255;255;255m$\033[0m                     \033[38;2;255;255;255m$$$$$$$$$$\033[0m                                             \033[0m");
  $display("\033[0m                                              \033[38;2;255;255;255m$$$\033[38;2;255;244;234mB\033[38;2;239;205;175ma\033[38;2;226;217;206m#\033[38;2;255;255;255m$\033[0m                   \033[38;2;255;255;255m$$$\033[38;2;255;251;252m$\033[38;2;255;227;227m8\033[38;2;255;215;212mW\033[38;2;255;207;200m#\033[38;2;255;203;188m*\033[38;2;255;203;178m*\033[38;2;255;228;208m&\033[38;2;255;255;255m$$$$\033[0m                                           \033[0m");
  $display("\033[0m                                         \033[38;2;255;255;255m$\033[38;2;248;255;255m$\033[38;2;238;240;240m%%\033[38;2;226;225;222mM\033[38;2;234;228;221mW\033[38;2;246;236;227m8\033[38;2;246;236;228m8\033[38;2;238;231;223m&\033[38;2;217;211;204mo\033[38;2;197;171;152mw\033[38;2;235;201;177ma\033[38;2;207;203;199ma\033[38;2;217;214;212m*\033[38;2;230;225;221mW\033[38;2;241;238;233m8\033[38;2;247;247;243mB\033[38;2;246;249;252m@\033[38;2;255;255;255m$$\033[0m          \033[38;2;255;255;255m$$$\033[38;2;255;252;254m$\033[38;2;251;165;172mk\033[38;2;247;143;148mq\033[38;2;250;184;182ma\033[38;2;248;160;143mp\033[38;2;247;159;129mq\033[38;2;251;204;185m*\033[38;2;252;217;198mM\033[38;2;245;141;58mL\033[38;2;247;160;71mO\033[38;2;255;245;230mB\033[38;2;255;255;255m$$\033[0m                                           \033[0m");
  $display("\033[0m                                      \033[38;2;255;255;255m$$\033[38;2;223;225;226mM\033[38;2;209;204;199ma\033[38;2;225;209;194mo\033[38;2;235;208;188mo\033[38;2;240;206;184mo\033[38;2;241;205;182mo\033[38;2;222;189;168mb\033[38;2;206;175;156mq\033[38;2;202;171;152mw\033[38;2;197;165;147mm\033[38;2;205;172;156mq\033[38;2;249;208;188m*\033[38;2;219;184;165mb\033[38;2;180;156;139mO\033[38;2;203;176;157mq\033[38;2;247;214;192m#\033[38;2;255;224;203mW\033[38;2;247;224;205mW\033[38;2;229;214;201m*\033[38;2;217;212;208m*\033[38;2;227;228;228mW\033[38;2;252;255;255m$\033[38;2;255;255;255m$\033[0m       \033[38;2;255;255;255m$$\033[38;2;255;249;249m@\033[38;2;245;112;119mO\033[38;2;244;99;100mL\033[38;2;254;245;246m@\033[38;2;251;197;180mo\033[38;2;242;95;39mX\033[38;2;243;110;38mY\033[38;2;253;228;213m&\033[38;2;255;255;255m$\033[38;2;248;183;105mq\033[38;2;244;135;0mY\033[38;2;251;217;162mo\033[38;2;255;255;255m$$$$$$$$\033[0m   \033[38;2;255;255;255m$$$$$$$\033[0m                           \033[0m");
  $display("\033[0m                                    \033[38;2;255;255;255m$\033[38;2;247;251;251m@\033[38;2;222;221;218m#\033[38;2;208;196;186mk\033[38;2;216;189;172mb\033[38;2;235;198;178ma\033[38;2;247;207;185m*\033[38;2;250;208;189m*\033[38;2;242;201;183mo\033[38;2;199;167;152mw\033[38;2;216;180;164md\033[38;2;237;196;179ma\033[38;2;247;204;186m*\033[38;2;249;206;189m*\033[38;2;250;207;189m*\033[38;2;247;206;187m*\033[38;2;250;208;190m#\033[38;2;245;203;186mo\033[38;2;214;178;163md\033[38;2;178;151;137m0\033[38;2;223;188;168mb\033[38;2;249;208;187m*\033[38;2;247;207;185m*\033[38;2;240;202;182mo\033[38;2;219;193;174mk\033[38;2;206;194;182mk\033[38;2;226;225;222mM\033[38;2;255;255;255m$$\033[0m     \033[38;2;255;255;255m$$\033[38;2;255;246;246m@\033[38;2;245;113;103m0\033[38;2;248;153;137mq\033[38;2;255;255;255m$\033[38;2;246;146;98mZ\033[38;2;243;109;24mX\033[38;2;247;156;84mZ\033[38;2;255;255;255m$\033[38;2;253;231;197mW\033[38;2;245;155;14mJ\033[38;2;247;176;48m0\033[38;2;255;247;230mB\033[38;2;255;255;255m$$$\033[38;2;255;254;244m@\033[38;2;255;252;229mB\033[38;2;255;251;237mB\033[38;2;255;255;253m$\033[38;2;255;255;255m$$$$$\033[38;2;253;253;250m$\033[38;2;248;251;240mB\033[38;2;251;255;243m@\033[38;2;250;253;245m@\033[38;2;255;255;255m$$$$\033[0m                         \033[0m");
  $display("\033[0m                            \033[38;2;255;255;255m$$$$$\033[38;2;246;246;246mB\033[38;2;232;234;234m&\033[38;2;218;217;210m*\033[38;2;204;199;189mk\033[38;2;221;205;188ma\033[38;2;232;200;178ma\033[38;2;245;204;183mo\033[38;2;251;207;188m*\033[38;2;248;206;188m*\033[38;2;247;206;187m*\033[38;2;248;206;187m*\033[38;2;246;203;185mo\033[38;2;247;204;186m*\033[38;2;250;206;189m*\033[38;2;248;205;188m*\033[38;2;247;204;188m*\033[38;2;246;204;188m**\033[38;2;247;205;188m*\033[38;2;244;201;185mo\033[38;2;240;198;183mo\033[38;2;251;209;193m#\033[38;2;235;196;180ma\033[38;2;213;177;163mp\033[38;2;248;206;189m*\033[38;2;250;208;189m*\033[38;2;251;208;190m#\033[38;2;251;207;188m*\033[38;2;245;204;182mo\033[38;2;227;197;174mh\033[38;2;195;183;172mp\033[38;2;194;190;187mb\033[38;2;225;225;225mW\033[38;2;240;240;240m%%\033[38;2;255;255;255m$$$$$$\033[38;2;255;249;248m@\033[38;2;254;241;237mB\033[38;2;253;234;222m8\033[38;2;244;126;40mJ\033[38;2;243;126;16mY\033[38;2;248;182;104mq\033[38;2;251;210;146mh\033[38;2;248;182;73mm\033[38;2;253;210;132mh\033[38;2;255;255;244m@\033[38;2;255;255;255m$$$\033[38;2;255;251;232mB\033[38;2;249;210;45mm\033[38;2;250;225;102mb\033[38;2;254;243;182mW\033[38;2;255;247;186mW\033[38;2;255;255;214m%%\033[38;2;255;255;252m$\033[38;2;255;255;231mB\033[38;2;242;251;182mW\033[38;2;228;244;156mo\033[38;2;224;242;165mo\033[38;2;222;242;177m*\033[38;2;177;228;118mw\033[38;2;147;220;96m0\033[38;2;151;225;128mm\033[38;2;230;251;227m8\033[38;2;255;255;255m$$$\033[0m                        \033[0m");
  $display("\033[0m                           \033[38;2;255;255;255m$\033[38;2;232;229;225mW\033[38;2;187;177;161mw\033[38;2;178;165;142mO\033[38;2;171;155;126mQ\033[38;2;154;137;105mU\033[38;2;147;134;102mY\033[38;2;153;142;106mU\033[38;2;180;151;117mQ\033[38;2;228;191;165mk\033[38;2;246;204;181mo\033[38;2;247;205;185m*\033[38;2;245;204;185mo\033[38;2;246;203;185mo\033[38;2;248;204;186m*\033[38;2;236;196;179ma\033[38;2;207;173;159mq\033[38;2;248;206;189m*\033[38;2;247;204;188m*\033[38;2;247;204;189m**\033[38;2;246;204;188m*\033[38;2;246;203;186mo\033[38;2;246;204;187m*\033[38;2;250;207;189m*\033[38;2;185;153;140mO\033[38;2;220;183;169mb\033[38;2;248;206;190m*\033[38;2;247;205;189m*\033[38;2;250;206;191m*\033[38;2;247;205;188m*\033[38;2;214;179;163md\033[38;2;230;191;175mh\033[38;2;250;207;190m*\033[38;2;246;203;187m*\033[38;2;249;209;190m#\033[38;2;242;210;188m*\033[38;2;193;159;132mO\033[38;2;168;145;114mC\033[38;2;143;130;107mY\033[38;2;155;134;109mU\033[38;2;178;159;133m0\033[38;2;184;169;147mZ\033[38;2;183;173;158mw\033[38;2;209;204;198ma\033[38;2;255;255;255m$$$\033[38;2;250;197;149mh\033[38;2;244;129;9mY\033[38;2;245;148;21mJ\033[38;2;252;228;192mM\033[38;2;254;243;224m%%\033[38;2;255;255;253m$\033[38;2;255;255;255m$$$$$\033[38;2;255;254;251m$\033[38;2;252;239;173mM\033[38;2;251;234;122mh\033[38;2;253;245;172mM\033[38;2;251;249;197m&\033[38;2;238;238;118mh\033[38;2;223;232;74mq\033[38;2;217;233;98mp\033[38;2;235;244;177m#\033[38;2;249;252;233mB\033[38;2;236;248;221m8\033[38;2;173;227;130mq\033[38;2;124;213;77mJ\033[38;2;120;214;96mC\033[38;2;185;234;179mh\033[38;2;252;255;251m$\033[38;2;255;255;255m$$$\033[0m                        \033[0m");
  $display("\033[0m                           \033[38;2;255;255;255m$\033[38;2;207;197;178mk\033[38;2;107;72;22m-\033[38;2;110;74;26m?\033[38;2;98;67;25m-\033[38;2;111;98;61mr\033[38;2;168;153;92mJ\033[38;2;186;168;136mZ\033[38;2;247;231;217m&\033[38;2;247;214;197m#\033[38;2;244;202;182mo\033[38;2;245;203;185mo\033[38;2;246;203;187m*\033[38;2;246;203;188m*\033[38;2;251;206;190m*\033[38;2;181;150;137m0\033[38;2;220;183;169mb\033[38;2;248;206;190m*\033[38;2;246;203;187m*\033[38;2;246;203;186mo\033[38;2;245;203;187mo\033[38;2;245;202;187mo\033[38;2;245;203;186mo\033[38;2;247;203;186m*\033[38;2;240;197;180ma\033[38;2;165;137;126mC\033[38;2;246;203;187m*\033[38;2;246;203;186moo\033[38;2;246;202;187mo\033[38;2;247;203;188m*\033[38;2;235;194;179mh\033[38;2;176;147;136m0\033[38;2;232;191;177mh\033[38;2;250;205;190m*\033[38;2;246;203;187m*\033[38;2;249;226;212mW\033[38;2;254;238;225m%%\033[38;2;208;177;154mq\033[38;2;174;144;93mJ\033[38;2;141;129;83mz\033[38;2;95;64;28m_\033[38;2;112;75;27m?\033[38;2;107;72;23m-\033[38;2;143;127;101mX\033[38;2;255;255;255m$$\033[38;2;255;253;250m$\033[38;2;246;163;61m0\033[38;2;244;141;0mY\033[38;2;248;182;67mZ\033[38;2;255;255;255m$$$$\033[0m  \033[38;2;255;255;255m$$$$\033[38;2;252;248;190m&\033[38;2;239;233;61mq\033[38;2;226;229;39mZ\033[38;2;224;234;97md\033[38;2;221;237;134mk\033[38;2;221;240;170mo\033[38;2;228;245;202mW\033[38;2;208;239;181mo\033[38;2;141;217;88mL\033[38;2;115;212;79mJ\033[38;2;149;224;137mm\033[38;2;228;247;228m8\033[38;2;255;255;255m$$$\033[0m                          \033[0m");
  $display("\033[0m                           \033[38;2;255;255;255m$\033[38;2;211;207;199ma\033[38;2;96;66;26m_\033[38;2;83;57;28m+\033[38;2;133;123;81mv\033[38;2;169;150;95mJ\033[38;2;199;181;155mq\033[38;2;254;241;230m%%\033[38;2;250;234;220m8\033[38;2;245;208;193m*\033[38;2;246;202;185mo\033[38;2;248;205;188m*\033[38;2;246;203;188m*\033[38;2;247;207;191m*\033[38;2;224;184;169mb\033[38;2;176;145;132mQ\033[38;2;250;207;190m*\033[38;2;246;203;186moo\033[38;2;246;203;185mo\033[38;2;245;202;186moo\033[38;2;246;202;185mo\033[38;2;249;205;188m*\033[38;2;221;182;166mb\033[38;2;177;148;137m0\033[38;2;251;207;191m#\033[38;2;246;203;186mo\033[38;2;246;203;185mo\033[38;2;247;202;186mo\033[38;2;246;201;185mo\033[38;2;249;203;188m*\033[38;2;233;190;176mh\033[38;2;172;143;132mQ\033[38;2;247;204;188m*\033[38;2;249;218;204mM\033[38;2;247;215;201mM\033[38;2;249;232;219m&\033[38;2;255;243;231mB\033[38;2;212;182;159mp\033[38;2;178;144;92mJ\033[38;2;133;123;82mv\033[38;2;87;59;28m+\033[38;2;99;67;30m-\033[38;2;189;182;172mp\033[38;2;255;255;255m$$\033[38;2;254;239;218m8\033[38;2;247;169;43m0\033[38;2;247;172;37mQ\033[38;2;252;223;164m*\033[38;2;255;255;255m$$$\033[0m  \033[38;2;255;255;255m$$$\033[38;2;254;250;207m8\033[38;2;245;237;87mb\033[38;2;230;228;26mO\033[38;2;229;235;94md\033[38;2;245;249;209m8\033[38;2;255;255;255m$$\033[38;2;224;244;197mM\033[38;2;152;220;92m0\033[38;2;120;212;74mJ\033[38;2;118;214;97mC\033[38;2;158;227;156mp\033[38;2;250;254;251m@\033[38;2;255;255;255m$$$\033[0m  \033[38;2;255;255;255m$$$$$\033[0m                    \033[0m");
  $display("\033[0m                  \033[38;2;255;255;255m$$\033[0m       \033[38;2;255;255;255m$\033[38;2;229;229;229mW\033[38;2;87;71;52m?\033[38;2;145;126;74mc\033[38;2;162;134;74mX\033[38;2;195;175;156mw\033[38;2;255;243;230m%%\033[38;2;252;239;225m8\033[38;2;251;235;222m8\033[38;2;245;211;195m#\033[38;2;242;200;185mo\033[38;2;219;181;169mb\033[38;2;247;215;203mM\033[38;2;252;228;215m&\033[38;2;189;158;144mZ\033[38;2;218;180;165md\033[38;2;250;205;188m*\033[38;2;247;203;185mo\033[38;2;246;203;186mo\033[38;2;246;203;185mo\033[38;2;246;203;186moo\033[38;2;247;202;186mo\033[38;2;250;205;189m*\033[38;2;213;177;162mp\033[38;2;178;148;136m0\033[38;2;252;206;188m*\033[38;2;246;202;185mo\033[38;2;248;203;186m*\033[38;2;249;204;187m*\033[38;2;246;201;186mo\033[38;2;246;205;191m*\033[38;2;251;218;205mM\033[38;2;203;167;154mw\033[38;2;192;161;147mZ\033[38;2;254;227;213m&\033[38;2;248;226;213mW\033[38;2;246;208;193m*\033[38;2;247;225;212mW\033[38;2;254;237;224m8\033[38;2;209;168;148mw\033[38;2;164;128;81mX\033[38;2;131;111;63mn\033[38;2;175;165;154mZ\033[38;2;255;255;255m$$$$\033[38;2;255;255;249m$\033[38;2;255;255;251m$\033[38;2;255;255;255m$$$\033[0m   \033[38;2;255;255;255m$$\033[38;2;252;249;195m&\033[38;2;237;230;30mZ\033[38;2;225;228;38mZ\033[38;2;238;243;165m*\033[38;2;254;255;254m$\033[38;2;255;255;255m$\033[38;2;252;254;249m@\033[38;2;206;238;177mo\033[38;2;140;218;91mQ\033[38;2;114;212;81mJ\033[38;2;151;224;140mw\033[38;2;230;248;230m8\033[38;2;249;253;250m@\033[38;2;255;255;255m$$$\033[0m \033[38;2;255;255;255m$$$\033[38;2;251;253;253m$\033[38;2;246;250;252m@\033[38;2;253;253;255m$\033[38;2;255;255;255m$$$$\033[0m                 \033[0m");
  $display("\033[0m               \033[38;2;255;255;255m$$\033[38;2;245;243;241mB\033[38;2;231;229;223mW\033[38;2;253;251;245m@\033[38;2;253;253;253m$\033[38;2;255;255;255m$\033[0m     \033[38;2;255;255;255m$$\033[38;2;140;138;132mJ\033[38;2;148;117;63mv\033[38;2;195;166;139mZ\033[38;2;252;236;223m8\033[38;2;245;219;203mM\033[38;2;247;222;207mW\033[38;2;244;210;195m#\033[38;2;249;204;188m*\033[38;2;182;154;141mO\033[38;2;217;182;166md\033[38;2;248;219;205mM\033[38;2;250;215;199mM\033[38;2;185;153;141mO\033[38;2;223;185;170mb\033[38;2;249;204;187m*\033[38;2;247;201;184mo\033[38;2;246;202;186mooo\033[38;2;246;201;185mo\033[38;2;247;201;185mo\033[38;2;248;203;187m*\033[38;2;225;184;168mb\033[38;2;163;135;124mC\033[38;2;252;206;188m*\033[38;2;248;203;185m*\033[38;2;229;188;173mk\033[38;2;223;183;168mb\033[38;2;251;205;189m*\033[38;2;246;202;188m*\033[38;2;246;209;194m#\033[38;2;250;204;188m*\033[38;2;170;141;130mL\033[38;2;230;190;174mh\033[38;2;238;198;181ma\033[38;2;211;174;160mp\033[38;2;248;205;187m*\033[38;2;246;207;191m*\033[38;2;249;206;190m*\033[38;2;214;168;146mq\033[38;2;159;117;71mc\033[38;2;215;209;193ma\033[38;2;255;255;255m$\033[0m \033[38;2;255;255;255m$$$$$$$$\033[38;2;243;243;246mB\033[38;2;255;255;255m$$$\033[38;2;251;250;213m8\033[38;2;229;235;98md\033[38;2;242;247;194mW\033[38;2;255;255;255m$$\033[38;2;252;255;249m$\033[38;2;184;231;147md\033[38;2;120;212;76mJ\033[38;2;121;215;101mL\033[38;2;193;237;190ma\033[38;2;253;255;254m$\033[38;2;255;255;255m$$$$$$$$\033[38;2;159;211;231mh\033[38;2;90;175;217mO\033[38;2;73;163;221mQ\033[38;2;93;171;229mZ\033[38;2;145;198;238mb\033[38;2;227;243;255m%%\033[38;2;255;255;255m$$$\033[0m                \033[0m");
  $display("\033[0m            \033[38;2;255;255;255m$$\033[38;2;240;240;237m%%\033[38;2;243;242;235m%%\033[38;2;229;226;217mM\033[38;2;253;249;236mB\033[38;2;170;166;156mZ\033[38;2;227;223;210m#\033[38;2;205;202;193mh\033[38;2;211;210;207mo\033[38;2;240;240;242m%%\033[38;2;255;255;255m$\033[0m    \033[38;2;255;255;255m$\033[38;2;203;203;201mh\033[38;2;165;129;102mU\033[38;2;251;211;192m#\033[38;2;246;205;189m*\033[38;2;242;198;183mo\033[38;2;231;190;175mh\033[38;2;251;205;189m*\033[38;2;203;168;154mw\033[38;2;183;153;140mO\033[38;2;228;188;172mk\033[38;2;246;200;183mo\033[38;2;250;203;186m*\033[38;2;212;173;157mp\033[38;2;177;147;135m0\033[38;2;252;206;189m*\033[38;2;246;201;185mo\033[38;2;247;201;187mo\033[38;2;247;201;186mo\033[38;2;246;201;186mo\033[38;2;246;201;185mo\033[38;2;249;203;186m*\033[38;2;250;204;186m*\033[38;2;240;196;179ma\033[38;2;150;124;114mY\033[38;2;246;201;184mo\033[38;2;248;202;185mo\033[38;2;240;197;181ma\033[38;2;146;121;112mY\033[38;2;227;186;170mk\033[38;2;250;204;186m*\033[38;2;246;201;183mo\033[38;2;250;204;186m*\033[38;2;220;181;165md\033[38;2;175;145;134mQ\033[38;2;246;201;184mo\033[38;2;175;146;133mQ\033[38;2;246;203;184mo\033[38;2;246;202;185mo\033[38;2;247;201;185mo\033[38;2;251;207;189m*\033[38;2;204;160;132mZ\033[38;2;226;219;208m#\033[38;2;255;255;255m$\033[0m     \033[38;2;255;255;255m$\033[38;2;238;238;238m8\033[38;2;215;215;214m*\033[38;2;212;209;202mo\033[38;2;199;197;189mk\033[38;2;185;183;178mp\033[38;2;241;239;235m8\033[38;2;249;249;249m@\033[38;2;255;255;255m$$$$$\033[38;2;255;255;253m$\033[38;2;254;255;250m$\033[38;2;226;252;221m&\033[38;2;241;255;240mB\033[38;2;255;255;255m$$$\033[38;2;210;239;229mW\033[38;2;151;215;200md\033[38;2;142;212;204md\033[38;2;185;230;231m*\033[38;2;253;255;255m$\033[38;2;255;255;255m$\033[38;2;171;214;234ma\033[38;2;42;149;208mU\033[38;2;43;146;217mJ\033[38;2;111;180;230mw\033[38;2;203;227;246mW\033[38;2;206;229;246mW\033[38;2;124;184;227mq\033[38;2;185;216;239m*\033[38;2;255;255;255m$$$\033[0m               \033[0m");
  $display("\033[0m            \033[38;2;255;255;255m$\033[38;2;242;241;240m%%\033[38;2;208;204;190mh\033[38;2;202;196;185mk\033[38;2;193;188;179md\033[38;2;164;161;155mO\033[38;2;172;167;160mZ\033[38;2;184;180;172mq\033[38;2;212;207;197ma\033[38;2;239;234;222m&\033[38;2;219;216;211m*\033[38;2;249;249;249m@\033[38;2;255;255;255m$\033[0m   \033[38;2;255;255;255m$\033[38;2;212;209;205mo\033[38;2;224;188;168mb\033[38;2;249;205;187m*\033[38;2;249;205;189m*\033[38;2;213;175;161mp\033[38;2;203;167;153mw\033[38;2;240;197;181ma\033[38;2;166;139;127mL\033[38;2;241;198;181ma\033[38;2;168;140;129mL\033[38;2;250;203;185m*\033[38;2;252;206;189m*\033[38;2;194;157;144mZ\033[38;2;122;98;90mn\033[38;2;236;195;179ma\033[38;2;251;204;189m*\033[38;2;247;201;187mo\033[38;2;246;201;187mo\033[38;2;246;200;189mo\033[38;2;249;202;190m*\033[38;2;208;171;158mq\033[38;2;223;183;167mb\033[38;2;255;209;192m#\033[38;2;163;132;121mJ\033[38;2;214;176;162mp\033[38;2;250;203;186m*\033[38;2;255;209;191m#\033[38;2;157;126;115mU\033[38;2;141;112;103mz\033[38;2;231;191;175mh\033[38;2;251;204;187m*\033[38;2;247;201;184mo\033[38;2;251;205;187m*\033[38;2;163;134;123mC\033[38;2;229;189;173mk\033[38;2;175;145;133mQ\033[38;2;237;194;177mh\033[38;2;247;203;185mo\033[38;2;241;198;182mo\033[38;2;233;190;176mh\033[38;2;242;201;181mo\033[38;2;236;227;220mW\033[38;2;255;255;255m$\033[0m   \033[38;2;255;255;255m$\033[38;2;253;253;253m$\033[38;2;193;192;190mb\033[38;2;213;210;201mo\033[38;2;200;196;187mk\033[38;2;206;200;191mh\033[38;2;173;169;162mm\033[38;2;202;195;186mk\033[38;2;218;211;199mo\033[38;2;200;196;188mk\033[38;2;235;234;229m&\033[38;2;251;251;252m@\033[38;2;255;255;255m$$$$$$$$$\033[38;2;189;230;219m*\033[38;2;65;182;155mU\033[38;2;113;198;186mZ\033[38;2;154;212;210mb\033[38;2;129;199;209mq\033[38;2;164;213;226mh\033[38;2;255;255;255m$\033[38;2;93;172;225mZ\033[38;2;43;144;218mJ\033[38;2;71;158;222mQ\033[38;2;245;250;253m@\033[38;2;222;237;247m8\033[38;2;182;214;238mo\033[38;2;96;166;216mO\033[38;2;111;174;219mm\033[38;2;255;255;255m$$$\033[0m               \033[0m");
  $display("\033[0m            \033[38;2;255;255;255m$\033[38;2;233;233;232m&\033[38;2;226;220;208m#\033[38;2;185;180;172mq\033[38;2;212;207;197ma\033[38;2;144;141;135mC\033[38;2;136;133;127mU\033[38;2;187;181;175mp\033[38;2;252;249;237mB\033[38;2;254;248;235mB\033[38;2;253;250;243m@\033[38;2;252;252;252m$\033[38;2;255;255;255m$\033[0m  \033[38;2;255;255;255m$\033[38;2;238;239;240m%%\033[38;2;205;184;167md\033[38;2;250;206;188m*\033[38;2;246;203;188m*\033[38;2;250;207;191m#\033[38;2;186;154;141mO\033[38;2;226;186;171mk\033[38;2;189;157;145mZ\033[38;2;210;173;161mp\033[38;2;245;201;186mo\033[38;2;136;119;111mX\033[38;2;190;161;149mZ\033[38;2;245;200;187mo\033[38;2;190;155;144mZ\033[38;2;190;179;170mq\033[38;2;186;168;159mw\033[38;2;224;184;172mb\033[38;2;249;202;190m*\033[38;2;251;204;192m*\033[38;2;248;202;190m*\033[38;2;249;204;191m*\033[38;2;218;179;166md\033[38;2;120;104;97mu\033[38;2;204;173;162mq\033[38;2;202;165;152mw\033[38;2;127;112;104mc\033[38;2;196;171;159mw\033[38;2;214;176;163mp\033[38;2;208;170;158mq\033[38;2;158;136;125mJ\033[38;2;171;147;136mQ\033[38;2;215;179;164md\033[38;2;252;205;189m*\033[38;2;254;207;189m#\033[38;2;188;155;142mO\033[38;2;206;170;156mq\033[38;2;185;153;141mO\033[38;2;229;188;172mk\033[38;2;251;205;188m*\033[38;2;214;175;160mp\033[38;2;196;162;149mm\033[38;2;251;206;189m*\033[38;2;198;179;171mp\033[38;2;246;248;250m@\033[38;2;255;255;255m$\033[0m  \033[38;2;255;255;255m$\033[38;2;226;226;226mW\033[38;2;184;179;170mq\033[38;2;255;253;241m@\033[38;2;241;235;225m&\033[38;2;177;172;166mw\033[38;2;190;186;178mp\033[38;2;129;126;120mX\033[38;2;184;179;171mq\033[38;2;217;210;199mo\033[38;2;192;186;174mp\033[38;2;237;235;229m&\033[38;2;255;255;255m$\033[0m      \033[38;2;255;255;255m$$\033[38;2;201;234;229mM\033[38;2;88;185;182mQ\033[38;2;245;251;252m@\033[38;2;255;255;255m$$\033[38;2;234;244;251mB\033[38;2;143;197;236mb\033[38;2;47;145;218mJ\033[38;2;37;139;213mY\033[38;2;123;184;228mq\033[38;2;255;255;255m$\033[38;2;225;241;252m%%\033[38;2;159;205;238mh\033[38;2;180;216;242m*\033[38;2;250;255;255m$\033[38;2;255;255;255m$$$\033[0m               \033[0m");
  $display("\033[0m            \033[38;2;255;255;255m$$\033[38;2;235;234;230m&\033[38;2;204;201;191mh\033[38;2;190;185;175mp\033[38;2;221;215;204m*\033[38;2;228;223;213mM\033[38;2;196;191;185mb\033[38;2;254;249;238mB\033[38;2;252;247;238mB\033[38;2;250;249;248m@\033[38;2;255;255;255m$\033[0m  \033[38;2;255;255;255m$$\033[38;2;181;177;174mq\033[38;2;222;184;164mb\033[38;2;252;207;191m#\033[38;2;245;202;187mo\033[38;2;248;204;189m*\033[38;2;176;145;133mQ\033[38;2;232;191;176mh\033[38;2;167;139;128mL\033[38;2;222;183;168mb\033[38;2;167;150;139mQ\033[38;2;182;176;167mw\033[38;2;181;179;175mq\033[38;2;191;180;176mp\033[38;2;180;164;157mm\033[38;2;173;170;166mm\033[38;2;206;204;198mh\033[38;2;195;187;180md\033[38;2;194;172;164mq\033[38;2;207;173;163mp\033[38;2;228;189;176mk\033[38;2;241;199;185mo\033[38;2;247;202;187m*\033[38;2;159;138;129mC\033[38;2;199;196;189mk\033[38;2;206;197;188mk\033[38;2;145;139;135mJ\033[38;2;187;184;179mp\033[38;2;183;180;179mp\033[38;2;195;189;188mb\033[38;2;181;177;175mq\033[38;2;185;179;175mq\033[38;2;142;133;128mU\033[38;2;182;155;146mO\033[38;2;241;198;183mo\033[38;2;226;185;171mk\033[38;2;184;152;141mO\033[38;2;180;151;140m0\033[38;2;232;191;175mh\033[38;2;253;206;188m*\033[38;2;189;156;142mZ\033[38;2;224;185;169mb\033[38;2;253;208;190m#\033[38;2;174;146;132mQ\033[38;2;229;221;215mM\033[38;2;255;255;255m$\033[0m  \033[38;2;255;255;255m$\033[38;2;235;235;235m8\033[38;2;231;226;217mM\033[38;2;255;249;238mB\033[38;2;248;244;234m%%\033[38;2;158;155;148m0\033[38;2;166;163;156mO\033[38;2;195;192;184mb\033[38;2;210;206;197ma\033[38;2;185;180;171mq\033[38;2;228;223;214mM\033[38;2;237;236;234m8\033[38;2;255;255;255m$\033[0m      \033[38;2;255;255;255m$$$\033[38;2;192;227;234m#\033[38;2;123;193;217mq\033[38;2;133;194;229md\033[38;2;115;183;231mq\033[38;2;69;157;223mQ\033[38;2;35;139;214mY\033[38;2;42;141;213mU\033[38;2;93;167;221mO\033[38;2;227;240;249m8\033[38;2;255;255;255m$$$$$$\033[0m                 \033[0m");
  $display("\033[0m              \033[38;2;255;255;255m$\033[38;2;252;252;250m@\033[38;2;254;250;243m@\033[38;2;255;249;240m@\033[38;2;245;239;230m8\033[38;2;216;211;204mo\033[38;2;220;215;208m*\033[38;2;255;250;242m@\033[38;2;255;255;255m$$\033[0m  \033[38;2;255;255;255m$\033[38;2;240;240;239m%%\033[38;2;150;133;121mU\033[38;2;240;198;181ma\033[38;2;217;179;165md\033[38;2;245;202;187mo\033[38;2;248;204;189m*\033[38;2;175;144;134mQ\033[38;2;217;179;166md\033[38;2;143;125;116mY\033[38;2;160;148;141mQ\033[38;2;178;177;175mq\033[38;2;234;234;234m8\033[38;2;218;218;219m#\033[38;2;182;183;184mp\033[38;2;251;252;252m@\033[38;2;244;244;244mB\033[38;2;213;213;212m*\033[38;2;180;178;176mq\033[38;2;213;209;203mo\033[38;2;226;220;212m#\033[38;2;200;189;181mb\033[38;2;194;176;168mq\033[38;2;197;176;168mp\033[38;2;178;163;155mZ\033[38;2;196;191;185mb\033[38;2;196;193;188mb\033[38;2;211;210;210mo\033[38;2;245;246;246mB\033[38;2;255;255;255m$$\033[38;2;230;231;231m&\033[38;2;156;156;157m0\033[38;2;227;227;228mW\033[38;2;162;162;162mZ\033[38;2;157;147;142mL\033[38;2;198;170;160mq\033[38;2;173;143;132mQ\033[38;2;178;148;138m0\033[38;2;239;195;180ma\033[38;2;236;193;178mh\033[38;2;183;151;139m0\033[38;2;247;203;186m*\033[38;2;251;207;189m*\033[38;2;184;153;139mO\033[38;2;219;190;174mk\033[38;2;251;246;243mB\033[38;2;255;255;255m$\033[0m \033[38;2;255;255;255m$\033[38;2;251;251;251m@\033[38;2;249;245;236mB\033[38;2;252;247;237mB\033[38;2;226;221;212m#\033[38;2;222;217;209m#\033[38;2;248;243;234m%%\033[38;2;217;213;204mo\033[38;2;182;179;170mq\033[38;2;201;197;187mk\033[38;2;232;232;231m&\033[38;2;255;255;255m$\033[0m        \033[38;2;255;255;255m$$$\033[38;2;243;254;255m@\033[38;2;174;216;243mo\033[38;2;127;188;233mp\033[38;2;119;183;230mq\033[38;2;142;194;232mb\033[38;2;194;222;242m#\033[38;2;251;253;254m$\033[38;2;255;255;255m$$$\033[0m                     \033[0m");
  $display("\033[0m               \033[38;2;255;255;255m$$\033[38;2;247;248;248mB\033[38;2;224;221;216m#\033[38;2;230;224;214mM\033[38;2;245;239;230m8\033[38;2;252;246;238mB\033[38;2;252;249;243m@\033[38;2;247;247;245mB\033[38;2;255;255;255m$\033[0m \033[38;2;255;255;255m$\033[38;2;239;230;220mW\033[38;2;166;140;123mC\033[38;2;251;206;189m*\033[38;2;173;143;133mQ\033[38;2;236;194;180ma\033[38;2;252;205;191m#\033[38;2;183;150;140m0\033[38;2;202;168;155mw\033[38;2;143;136;131mJ\033[38;2;191;190;188mb\033[38;2;251;251;251m@\033[38;2;255;255;255m$\033[38;2;188;187;188md\033[38;2;112;112;112mv\033[38;2;252;252;252m$\033[38;2;255;255;255m$$\033[38;2;247;247;247mB\033[38;2;160;158;157mO\033[38;2;241;236;227m8\033[38;2;255;253;243m@\033[38;2;255;249;240m@\033[38;2;252;247;237mB\033[38;2;255;253;244m@\033[38;2;203;198;194mh\033[38;2;210;209;210mo\033[38;2;255;255;255m$$$$\033[38;2;208;208;208mo\033[38;2;107;107;107mu\033[38;2;245;245;245mB\033[38;2;255;255;255m$\033[38;2;173;173;173mw\033[38;2;194;189;183md\033[38;2;170;148;139mQ\033[38;2;180;148;137m0\033[38;2;249;203;188m*\033[38;2;185;153;142mO\033[38;2;222;183;168mb\033[38;2;249;205;187m*\033[38;2;252;207;190m#\033[38;2;178;148;137m0\033[38;2;215;178;162md\033[38;2;247;223;210mW\033[38;2;255;255;255m$$\033[38;2;250;248;248m@\033[38;2;249;246;240mB\033[38;2;252;247;237mB\033[38;2;246;241;232m%%\033[38;2;190;186;180md\033[38;2;211;206;199ma\033[38;2;227;222;215mM\033[38;2;234;230;223mW\033[38;2;225;222;218mM\033[38;2;240;240;238m%%\033[38;2;255;255;255m$\033[0m          \033[38;2;255;255;255m$$$$$$$\033[38;2;254;254;255m$\033[38;2;248;251;253m@\033[38;2;255;255;255m$$$$$$$$$$$\033[0m             \033[0m");
  $display("\033[0m                 \033[38;2;255;255;255m$\033[38;2;228;227;226mW\033[38;2;228;222;211m#\033[38;2;255;249;240m@\033[38;2;251;246;237mB\033[38;2;252;246;237mB\033[38;2;231;227;221mW\033[38;2;218;218;218m#\033[38;2;255;255;255m$\033[38;2;247;247;246mB\033[38;2;217;195;176mk\033[38;2;177;146;132mQ\033[38;2;255;208;193m#\033[38;2;205;168;156mq\033[38;2;196;162;150mm\033[38;2;255;210;194m#\033[38;2;194;159;150mm\033[38;2;178;149;138m0\033[38;2;127;123;119mX\033[38;2;247;247;248mB\033[38;2;255;255;255m$$$$$$$$\033[38;2;205;204;205ma\033[38;2;193;189;183md\033[38;2;255;253;243m@\033[38;2;252;247;237mBB\033[38;2;246;241;232m%%\033[38;2;179;177;175mq\033[38;2;255;255;255m$$$$$$$$$\033[38;2;217;216;217m#\033[38;2;177;174;169mw\033[38;2;164;148;138mQ\033[38;2;188;157;144mZ\033[38;2;218;181;167md\033[38;2;186;155;143mO\033[38;2;250;204;187m*\033[38;2;247;201;183mo\033[38;2;252;206;188m*\033[38;2;162;134;125mC\033[38;2;221;182;168mb\033[38;2;253;211;196m#\033[38;2;205;192;186mk\033[38;2;216;215;212m*\033[38;2;252;247;238mB\033[38;2;252;246;236mB\033[38;2;251;246;237mB\033[38;2;252;247;238mB\033[38;2;252;246;238mB\033[38;2;224;220;212m#\033[38;2;217;216;215m#\033[38;2;241;241;244m%%\033[38;2;255;255;255m$$\033[0m              \033[38;2;255;255;255m$$\033[38;2;222;237;247m8\033[38;2;106;171;217mZ\033[38;2;73;152;208mL\033[38;2;70;149;205mC\033[38;2;105;168;212mO\033[38;2;230;242;251m%%\033[38;2;255;255;255m$$\033[38;2;245;250;255m@\033[38;2;190;205;235mo\033[38;2;171;184;225mb\033[38;2;195;198;233mo\033[38;2;245;245;255m@\033[38;2;255;255;255m$$$\033[0m            \033[0m");
  $display("\033[0m                 \033[38;2;255;255;255m$\033[38;2;253;253;253m$\033[38;2;237;235;231m8\033[38;2;250;243;234m%%\033[38;2;252;246;238mBB\033[38;2;251;247;238mB\033[38;2;189;186;179mp\033[38;2;209;210;210mo\033[38;2;189;180;176mp\033[38;2;201;168;152mw\033[38;2;191;156;145mZ\033[38;2;252;206;191m#\033[38;2;244;199;185mo\033[38;2;167;140;130mL\033[38;2;244;199;184mo\033[38;2;226;185;171mk\033[38;2;139;118;110mX\033[38;2;131;127;123mY\033[38;2;252;252;252m$\033[38;2;255;255;255m$$$$$$$$\033[38;2;220;219;220m#\033[38;2;185;182;175mp\033[38;2;255;255;244m@\033[38;2;252;249;238mB\033[38;2;253;250;239mB\033[38;2;243;239;230m8\033[38;2;179;177;176mq\033[38;2;255;255;255m$$$$$$$$$\033[38;2;219;219;220m#\033[38;2;176;173;169mw\033[38;2;122;111;105mv\033[38;2;220;182;167mb\033[38;2;169;142;131mL\033[38;2;244;200;183mo\033[38;2;248;202;185mo\033[38;2;246;201;184mo\033[38;2;251;206;190m*\033[38;2;156;127;118mU\033[38;2;228;181;165mb\033[38;2;223;186;172mb\033[38;2;175;163;154mZ\033[38;2;238;233;224m&\033[38;2;253;248;238mB\033[38;2;252;246;237mBBB\033[38;2;249;244;238mB\033[38;2;243;243;243mB\033[38;2;255;255;255m$\033[0m                \033[38;2;255;255;255m$$$\033[38;2;110;173;218mm\033[38;2;120;179;221mw\033[38;2;203;225;241mM\033[38;2;201;224;240mM\033[38;2;105;167;210mO\033[38;2;148;191;222md\033[38;2;255;255;255m$\033[38;2;188;204;230mo\033[38;2;87;120;190mU\033[38;2;66;90;178mv\033[38;2;84;92;180mz\033[38;2;106;101;185mY\033[38;2;124;103;188mJ\033[38;2;207;193;229mo\033[38;2;255;255;255m$$$\033[0m           \033[0m");
  $display("\033[0m                  \033[38;2;255;255;255m$\033[38;2;250;250;251m@\033[38;2;235;231;225m&\033[38;2;252;246;238mB\033[38;2;252;246;237mB\033[38;2;252;247;238mB\033[38;2;255;251;241m@\033[38;2;191;187;181md\033[38;2;149;133;125mJ\033[38;2;197;165;152mw\033[38;2;209;172;159mp\033[38;2;250;204;188m**\033[38;2;214;175;163mp\033[38;2;181;150;140m0\033[38;2;255;209;195m#\033[38;2;147;124;117mY\033[38;2;122;121;116mz\033[38;2;229;228;229mW\033[38;2;255;255;255m$$$$$$$$\033[38;2;189;188;188md\033[38;2;215;210;203mo\033[38;2;255;253;241m@\033[38;2;255;252;240m@\033[38;2;253;250;238mB\033[38;2;254;252;240m@\033[38;2;185;182;177mp\033[38;2;221;221;222mM\033[38;2;255;255;255m$$$$$$$$\033[38;2;191;190;190mb\033[38;2;181;176;169mw\033[38;2;162;138;129mC\033[38;2;182;151;138m0\033[38;2;213;175;162mp\033[38;2;250;205;187m*\033[38;2;246;201;185mo\033[38;2;247;201;188m*\033[38;2;253;205;192m#\033[38;2;161;129;119mJ\033[38;2;178;135;118mC\033[38;2;188;179;171mq\033[38;2;248;244;235m%%\033[38;2;255;249;239mB\033[38;2;252;246;237mBBB\033[38;2;252;248;240mB\033[38;2;250;250;249m@\033[38;2;255;255;255m$\033[0m                 \033[38;2;255;255;255m$$$\033[38;2;122;178;218mw\033[38;2;163;202;230mh\033[38;2;253;255;253m$\033[38;2;255;255;255m$\033[38;2;243;247;251mB\033[38;2;204;218;237m#\033[38;2;138;163;210mm\033[38;2;70;101;182mz\033[38;2;76;90;178mc\033[38;2;146;148;206mZ\033[38;2;226;225;242m&\033[38;2;251;252;253m$\033[38;2;235;230;244m8\033[38;2;156;109;193mQ\033[38;2;243;235;247m%%\033[38;2;255;255;255m$$\033[0m           \033[0m");
  $display("\033[0m                   \033[38;2;255;255;255m$\033[38;2;224;224;223mM\033[38;2;226;221;211m#\033[38;2;255;249;239mB\033[38;2;252;245;236mB\033[38;2;253;245;236mB\033[38;2;255;251;242m@\033[38;2;206;198;190mh\033[38;2;132;114;108mz\033[38;2;230;188;174mk\033[38;2;247;201;187mo\033[38;2;244;199;185mo\033[38;2;250;204;190m*\033[38;2;203;168;157mq\033[38;2;189;157;147mZ\033[38;2;219;180;168mb\033[38;2;151;145;140mL\033[38;2;180;179;178mq\033[38;2;244;243;244mB\033[38;2;255;255;255m$$$$$\033[38;2;251;251;252m@\033[38;2;213;213;213m*\033[38;2;182;180;176mq\033[38;2;252;249;239mB\033[38;2;253;249;238mB\033[38;2;224;220;211m#\033[38;2;251;247;236mB\033[38;2;253;250;238mB\033[38;2;246;243;234m%%\033[38;2;185;183;180mp\033[38;2;201;200;199mh\033[38;2;237;237;237m8\033[38;2;252;252;252m$\033[38;2;255;255;255m$$\033[38;2;251;251;252m@\033[38;2;233;232;233m&\033[38;2;200;199;198mh\033[38;2;189;186;181md\033[38;2;160;144;136mL\033[38;2;173;142;131mL\033[38;2;188;154;144mZ\033[38;2;252;206;189m*\033[38;2;245;200;183mo\033[38;2;244;199;184mo\033[38;2;246;200;189mo\033[38;2;252;204;193m#\033[38;2;154;129;122mJ\033[38;2;196;188;180md\033[38;2;255;250;241m@\033[38;2;255;247;237mB\033[38;2;253;246;236mB\033[38;2;253;246;237mB\033[38;2;255;248;240mB\033[38;2;247;242;234m%%\033[38;2;249;249;247m@\033[38;2;255;255;255m$\033[0m                  \033[38;2;255;255;255m$$$\033[38;2;224;237;246m8\033[38;2;72;146;199mJ\033[38;2;67;137;196mU\033[38;2;87;140;199mC\033[38;2;83;126;192mU\033[38;2;69;104;183mz\033[38;2;66;89;177mv\033[38;2;94;100;184mY\033[38;2;179;177;220mb\033[38;2;255;255;255m$\033[38;2;207;190;227mo\033[38;2;187;155;212mp\033[38;2;192;150;211mp\033[38;2;166;102;191m0\033[38;2;245;237;248mB\033[38;2;255;255;255m$$\033[0m           \033[0m");
  $display("\033[0m                   \033[38;2;255;255;255m$\033[38;2;253;253;253m$\033[38;2;230;228;224mW\033[38;2;248;240;230m%%\033[38;2;254;246;237mB\033[38;2;255;248;238mB\033[38;2;251;246;237mB\033[38;2;167;152;145m0\033[38;2;115;85;77mr\033[38;2;237;195;180ma\033[38;2;244;199;184moo\033[38;2;245;200;186mo\033[38;2;250;204;190m*\033[38;2;203;167;156mw\033[38;2;188;157;146mZ\033[38;2;176;159;149mO\033[38;2;221;216;209m*\033[38;2;187;184;181mp\033[38;2;201;200;199mh\033[38;2;216;215;215m*\033[38;2;222;222;221mM\033[38;2;221;220;220m#\033[38;2;209;208;207mo\033[38;2;194;192;190mb\033[38;2;216;212;206mo\033[38;2;253;249;239mB\033[38;2;253;250;239mB\033[38;2;253;249;238mB\033[38;2;233;230;219mW\033[38;2;251;248;236mB\033[38;2;252;249;237mB\033[38;2;253;249;238mB\033[38;2;255;251;241m@\033[38;2;230;225;218mM\033[38;2;197;193;188mb\033[38;2;197;194;191mk\033[38;2;199;197;195mk\033[38;2;202;200;198mh\033[38;2;201;198;195mh\033[38;2;212;207;203mo\033[38;2;232;227;221mW\033[38;2;160;150;143mQ\033[38;2;146;122;114mY\033[38;2;189;156;145mZ\033[38;2;250;204;188m*\033[38;2;245;201;183mo\033[38;2;244;199;182mo\033[38;2;244;199;185mo\033[38;2;246;200;188mo\033[38;2;242;196;183mo\033[38;2;165;143;134mL\033[38;2;255;248;239mB\033[38;2;255;246;236mB\033[38;2;254;246;236mB\033[38;2;253;247;237mB\033[38;2;255;249;240m@\033[38;2;215;210;205mo\033[38;2;238;238;235m8\033[38;2;255;255;255m$\033[0m                    \033[38;2;255;255;255m$$$\033[38;2;246;253;255m@\033[38;2;169;198;229mh\033[38;2;128;160;210mZ\033[38;2;125;148;206mO\033[38;2;145;156;210mm\033[38;2;182;184;225mk\033[38;2;238;237;251m%%\033[38;2;255;255;255m$$\033[38;2;251;245;255m@\033[38;2;219;194;235m#\033[38;2;222;193;235m#\033[38;2;252;242;255m@\033[38;2;255;255;255m$$$\033[0m           \033[0m");
  $display("\033[0m                    \033[38;2;255;255;255m$\033[38;2;249;249;251m@\033[38;2;232;229;224mW\033[38;2;254;246;234mB\033[38;2;242;237;228m8\033[38;2;145;131;121mU\033[38;2;119;74;58mf\033[38;2;124;85;72mr\033[38;2;236;191;176mh\033[38;2;244;199;184mo\033[38;2;246;201;184mo\033[38;2;245;200;185mo\033[38;2;244;199;185mo\033[38;2;250;204;190m*\033[38;2;212;175;164mp\033[38;2;141;122;113mX\033[38;2;194;189;181md\033[38;2;255;254;243m@\033[38;2;238;232;223m&\033[38;2;231;225;216mM\033[38;2;228;222;215mM\033[38;2;230;224;217mM\033[38;2;239;233;225m&\033[38;2;249;244;235m%%\033[38;2;225;221;213m#\033[38;2;242;236;227m8\033[38;2;252;247;237mB\033[38;2;255;250;239m@\033[38;2;255;254;242m@\033[38;2;255;252;241m@@\033[38;2;253;249;238mB\033[38;2;244;239;230m8\033[38;2;221;216;209m*\033[38;2;248;242;233m%%\033[38;2;254;248;239mB\033[38;2;247;238;230m8\033[38;2;249;241;232m%%\033[38;2;255;247;237mB\033[38;2;249;244;235m%%\033[38;2;159;151;144mQ\033[38;2;153;130;121mU\033[38;2;223;184;171mb\033[38;2;251;205;190m*\033[38;2;245;200;185mo\033[38;2;244;200;184mo\033[38;2;245;200;184mo\033[38;2;246;201;184mo\033[38;2;246;202;186mo\033[38;2;230;177;160mb\033[38;2;169;150;140m0\033[38;2;255;250;239m@\033[38;2;254;246;236mB\033[38;2;255;247;237mB\033[38;2;255;250;240m@\033[38;2;194;185;177md\033[38;2;182;171;163mw\033[38;2;252;252;252m$\033[38;2;255;255;255m$\033[0m                     \033[38;2;255;255;255m$$$$$$$$$$$$$$$$$\033[0m            \033[0m");
  $display("\033[0m                     \033[38;2;255;255;255m$\033[38;2;240;240;240m%%\033[38;2;204;202;196mh\033[38;2;137;126;117mY\033[38;2;111;76;58mf\033[38;2;121;79;60mj\033[38;2;106;71;58mt\033[38;2;223;173;156mp\033[38;2;245;201;184mo\033[38;2;245;200;183mo\033[38;2;245;200;185mo\033[38;2;244;200;184moo\033[38;2;248;203;188m*\033[38;2;228;186;173mk\033[38;2;135;119;112mX\033[38;2;214;210;201mo\033[38;2;255;253;242m@\033[38;2;254;246;236mB\033[38;2;255;248;238mB\033[38;2;255;248;239mB\033[38;2;253;248;239mB\033[38;2;251;246;237mB\033[38;2;209;205;198ma\033[38;2;194;190;183mb\033[38;2;200;196;189mk\033[38;2;204;200;193mh\033[38;2;205;201;193mh\033[38;2;207;202;195mh\033[38;2;203;199;192mh\033[38;2;206;203;195mh\033[38;2;207;203;196mh\033[38;2;218;213;206m*\033[38;2;249;244;235m%%\033[38;2;252;246;237mB\033[38;2;253;245;235mB\033[38;2;255;247;237mB\033[38;2;248;243;233m%%\033[38;2;179;167;159mm\033[38;2;197;164;153mw\033[38;2;241;197;185mo\033[38;2;248;203;188m*\033[38;2;244;199;184mo\033[38;2;243;199;184mo\033[38;2;243;198;184mo\033[38;2;244;198;184mo\033[38;2;246;200;185mo\033[38;2;245;196;180mo\033[38;2;206;140;122m0\033[38;2;142;130;122mU\033[38;2;255;250;238mB\033[38;2;255;247;237mB\033[38;2;251;246;237mB\033[38;2;174;167;160mm\033[38;2;204;170;157mq\033[38;2;247;210;193m#\033[38;2;244;240;237m%%\033[38;2;255;255;255m$\033[0m                        \033[38;2;255;255;255m$$$$$\033[0m                     \033[0m");
  $display("\033[0m                      \033[38;2;255;255;255m$\033[38;2;163;159;156mO\033[38;2;102;73;56mt\033[38;2;113;80;61mf\033[38;2;110;75;58mf\033[38;2;97;65;52m?\033[38;2;188;133;115mL\033[38;2;247;200;181mo\033[38;2;243;198;183mo\033[38;2;244;199;184mo\033[38;2;246;201;184mo\033[38;2;246;201;185mo\033[38;2;244;199;185mo\033[38;2;247;202;188m*\033[38;2;242;198;184mo\033[38;2;180;158;150mZ\033[38;2;216;213;206mo\033[38;2;255;252;243m@\033[38;2;255;246;236mB\033[38;2;254;247;237mB\033[38;2;253;247;238mB\033[38;2;252;246;237mB\033[38;2;255;250;241m@\033[38;2;255;249;240m@\033[38;2;251;246;237mB\033[38;2;247;243;234m%%\033[38;2;243;239;230m8\033[38;2;240;236;227m8\033[38;2;244;239;230m8\033[38;2;250;245;236mB\033[38;2;254;248;239mB\033[38;2;255;249;240m@\033[38;2;252;246;238mB\033[38;2;251;246;237mB\033[38;2;253;247;238mB\033[38;2;252;248;239mB\033[38;2;178;169;162mm\033[38;2;218;180;168md\033[38;2;253;206;192m#\033[38;2;245;200;186mo\033[38;2;243;198;184moo\033[38;2;243;198;183moo\033[38;2;244;199;184mo\033[38;2;243;196;183mo\033[38;2;234;162;144mp\033[38;2;155;97;83mv\033[38;2;105;70;61mt\033[38;2;213;205;195ma\033[38;2;244;239;230m8\033[38;2;137;120;112mX\033[38;2;92;67;58m1\033[38;2;232;191;176mh\033[38;2;246;205;189m*\033[38;2;244;237;234m8\033[38;2;255;255;255m$\033[0m                                                  \033[0m");
  $display("\033[0m                     \033[38;2;255;255;255m$\033[38;2;216;215;214m*\033[38;2;112;91;74mr\033[38;2;108;79;61mf\033[38;2;99;71;57m1\033[38;2;99;70;56m1\033[38;2;98;66;53m1\033[38;2;136;86;74mx\033[38;2;240;173;154mb\033[38;2;246;199;184mo\033[38;2;244;198;183mo\033[38;2;244;200;184mo\033[38;2;245;201;185mo\033[38;2;245;200;186mo\033[38;2;243;199;185mo\033[38;2;245;200;187mo\033[38;2;246;200;189mo\033[38;2;187;159;152mZ\033[38;2;205;199;193mh\033[38;2;255;253;243m@\033[38;2;255;248;238mB\033[38;2;255;247;237mB\033[38;2;253;247;237mB\033[38;2;252;246;237mBBB\033[38;2;251;246;237mB\033[38;2;252;247;238mB\033[38;2;253;247;238mB\033[38;2;252;247;238mB\033[38;2;251;246;237mB\033[38;2;252;246;237mBB\033[38;2;253;246;238mB\033[38;2;254;248;238mB\033[38;2;255;252;242m@\033[38;2;191;184;176mp\033[38;2;206;172;161mq\033[38;2;250;204;191m*\033[38;2;244;199;185mo\033[38;2;243;199;184mo\033[38;2;243;198;184mo\033[38;2;243;198;183moo\033[38;2;243;199;184mo\033[38;2;243;195;181ma\033[38;2;234;160;145mq\033[38;2;185;111;100mU\033[38;2;104;62;51m1\033[38;2;112;67;53mt\033[38;2;113;98;91mn\033[38;2;116;105;96mu\033[38;2;86;52;35m+\033[38;2;87;56;43m_\033[38;2;205;167;154mw\033[38;2;224;191;176mk\033[38;2;233;232;231m&\033[38;2;255;255;255m$\033[0m                                                  \033[0m");
  $display("\033[0m                    \033[38;2;255;255;255m$\033[38;2;250;250;251m@\033[38;2;146;135;125mJ\033[38;2;105;79;62mf\033[38;2;97;73;60m1\033[38;2;90;66;55m?\033[38;2;91;65;53m?\033[38;2;100;68;56m1\033[38;2;93;60;51m?\033[38;2;182;113;99mU\033[38;2;243;180;163mk\033[38;2;246;199;184mo\033[38;2;243;198;183moo\033[38;2;244;200;184mo\033[38;2;244;199;184mo\033[38;2;244;199;185mo\033[38;2;244;200;186mo\033[38;2;249;202;190m*\033[38;2;178;152;143m0\033[38;2;202;197;189mk\033[38;2;246;241;231m%%\033[38;2;251;245;235mB\033[38;2;254;248;239mB\033[38;2;255;251;241m@\033[38;2;255;253;243m@\033[38;2;255;252;242m@@@\033[38;2;255;251;241m@\033[38;2;255;252;242m@@@@\033[38;2;255;251;241m@\033[38;2;250;246;236mB\033[38;2;209;205;197ma\033[38;2;184;156;146mZ\033[38;2;252;205;191m#\033[38;2;244;199;185mo\033[38;2;243;198;184mo\033[38;2;244;198;184mo\033[38;2;245;198;183mo\033[38;2;244;198;183mo\033[38;2;244;200;185mo\033[38;2;241;190;176mh\033[38;2;233;153;139mw\033[38;2;181;108;97mY\033[38;2;102;61;57m1\033[38;2;99;62;52m?\033[38;2;95;63;53m?\033[38;2;85;57;48m-\033[38;2;58;40;32m!\033[38;2;74;47;34m~\033[38;2;80;53;39m+\033[38;2;137;118;110mz\033[38;2;217;209;206mo\033[38;2;253;255;255m$\033[38;2;255;255;255m$\033[0m                                                  \033[0m");
  $display("\033[0m                    \033[38;2;255;255;255m$\033[38;2;218;215;212m*\033[38;2;110;89;72mr\033[38;2;102;78;65mf\033[38;2;93;69;58m1\033[38;2;88;64;53m?\033[38;2;89;62;51m-\033[38;2;91;63;52m?\033[38;2;95;64;54m?\033[38;2;104;68;59mt\033[38;2;208;128;112mQ\033[38;2;240;173;157mb\033[38;2;244;197;182mo\033[38;2;244;199;184mo\033[38;2;243;199;183moo\033[38;2;244;199;184mo\033[38;2;243;199;184mo\033[38;2;246;199;185mo\033[38;2;245;198;184mo\033[38;2;155;130;121mJ\033[38;2;142;112;101mz\033[38;2;166;133;122mC\033[38;2;172;143;131mL\033[38;2;163;144;135mL\033[38;2;168;155;147m0\033[38;2;198;182;172mp\033[38;2;198;183;171mp\033[38;2;201;187;176md\033[38;2;205;192;182mb\033[38;2;198;183;172mp\033[38;2;194;178;167mq\033[38;2;189;177;167mq\033[38;2;184;165;155mm\033[38;2;165;145;136mL\033[38;2;175;138;126mL\033[38;2;134;106;96mv\033[38;2;228;188;174mk\033[38;2;247;201;187mo\033[38;2;243;198;183mo\033[38;2;243;199;183moo\033[38;2;245;199;184mo\033[38;2;246;197;181mo\033[38;2;240;176;161mb\033[38;2;215;134;120m0\033[38;2;153;91;81mv\033[38;2;97;59;52m?\033[38;2;95;60;51m?\033[38;2;89;60;51m-\033[38;2;86;59;51m-\033[38;2;88;61;50m-\033[38;2;79;57;48m_\033[38;2;62;45;37mi\033[38;2;76;57;40m+\033[38;2;163;162;158mO\033[38;2;255;255;255m$\033[0m                                                    \033[0m");
  $display("\033[0m                    \033[38;2;255;255;255m$\033[38;2;200;193;184mb\033[38;2;105;82;60mf\033[38;2;101;79;64mf\033[38;2;92;69;57m1\033[38;2;88;64;53m?\033[38;2;87;63;53m-\033[38;2;86;61;50m-\033[38;2;90;63;50m-\033[38;2;91;61;50m-\033[38;2;109;70;63mt\033[38;2;197;116;105mJ\033[38;2;234;155;139mq\033[38;2;241;185;168mh\033[38;2;244;197;181mo\033[38;2;245;198;183mo\033[38;2;243;198;182mo\033[38;2;243;197;182moo\033[38;2;245;198;183mo\033[38;2;241;194;182ma\033[38;2;133;94;83mn\033[38;2;124;67;53mf\033[38;2;135;117;109mz\033[38;2;188;174;162mw\033[38;2;155;135;122mJ\033[38;2;209;168;145mw\033[38;2;197;155;132mO\033[38;2;195;155;132mO\033[38;2;195;156;133mO\033[38;2;199;158;136mZ\033[38;2;215;177;155mp\033[38;2;185;162;145mZ\033[38;2;180;163;153mZ\033[38;2;198;183;175md\033[38;2;103;85;81mj\033[38;2;145;115;106mX\033[38;2;251;205;189m*\033[38;2;244;198;184mo\033[38;2;245;198;184mo\033[38;2;245;199;184mo\033[38;2;245;197;183mo\033[38;2;243;181;168mk\033[38;2;220;144;132mZ\033[38;2;158;94;86mv\033[38;2;108;66;59mt\033[38;2;89;56;50m-\033[38;2;90;60;51m-\033[38;2;85;59;49m-\033[38;2;84;59;50m-\033[38;2;85;62;52m-\033[38;2;85;63;52m-\033[38;2;88;67;56m?\033[38;2;77;61;53m-\033[38;2;65;53;41m~\033[38;2;157;153;147mQ\033[38;2;255;255;255m$\033[0m                                                    \033[0m");
  $display("\033[0m                    \033[38;2;255;255;255m$\033[38;2;234;234;233m&\033[38;2;146;138;129mJ\033[38;2;96;77;61mt\033[38;2;95;75;59m1\033[38;2;88;67;55m?\033[38;2;84;60;49m-\033[38;2;89;62;52m-\033[38;2;87;60;49m-\033[38;2;87;61;50m-\033[38;2;87;60;50m-\033[38;2;94;62;55m?\033[38;2;142;86;77mn\033[38;2;188;114;100mU\033[38;2;229;151;133mw\033[38;2;242;177;160mb\033[38;2;246;192;176ma\033[38;2;247;197;182mo\033[38;2;245;197;181moo\033[38;2;250;201;186m*\033[38;2;196;158;146mZ\033[38;2;113;66;55mt\033[38;2;135;124;118mX\033[38;2;191;189;182md\033[38;2;178;171;163mm\033[38;2;226;206;190mo\033[38;2;246;219;199mM\033[38;2;243;216;197m#\033[38;2;246;220;202mM\033[38;2;246;226;212mW\033[38;2;226;215;204m*\033[38;2;204;197;188mk\033[38;2;206;202;193mh\033[38;2;158;154;148m0\033[38;2;94;60;52m?\033[38;2;170;134;124mC\033[38;2;253;203;188m*\033[38;2;248;199;185mo\033[38;2;247;194;180mo\033[38;2;239;175;159mb\033[38;2;213;140;127mO\033[38;2;162;99;90mz\033[38;2;109;66;60mt\033[38;2;90;57;50m-\033[38;2;88;58;49m-\033[38;2;85;58;51m-\033[38;2;82;58;51m-\033[38;2;81;59;51m-\033[38;2;83;61;50m-\033[38;2;85;64;53m-\033[38;2;85;65;54m?\033[38;2;89;69;56m?\033[38;2;98;79;63mt\033[38;2;86;70;53m?\033[38;2;137;133;125mU\033[38;2;255;255;255m$\033[0m                                                    \033[0m");
  $display("\033[0m                     \033[38;2;255;255;255m$$\033[38;2;187;185;183md\033[38;2;114;103;95mu\033[38;2;90;71;57m1\033[38;2;85;65;52m-\033[38;2;79;56;45m_\033[38;2;87;62;51m-\033[38;2;88;61;50m--\033[38;2;89;61;50m-\033[38;2;88;58;50m-\033[38;2;89;58;52m-\033[38;2;121;76;67mj\033[38;2;159;96;85mc\033[38;2;186;116;103mJ\033[38;2;211;141;129mO\033[38;2;230;163;148mp\033[38;2;241;179;163mk\033[38;2;251;191;176ma\033[38;2;221;175;164md\033[38;2;109;71;62mt\033[38;2;114;90;81mx\033[38;2;224;218;209m#\033[38;2;251;244;233m%%\033[38;2;251;243;233m%%\033[38;2;255;250;239m@@\033[38;2;255;251;240m@\033[38;2;255;249;238mB\033[38;2;241;235;224m&\033[38;2;252;245;234mB\033[38;2;239;233;223m&\033[38;2;112;93;85mx\033[38;2;110;69;55mt\033[38;2;141;110;102mz\033[38;2;232;175;163mb\033[38;2;205;145;133mO\033[38;2;177;115;104mU\033[38;2;135;83;75mx\033[38;2;93;59;54m?\033[38;2;76;51;47m+\033[38;2;86;57;51m-\033[38;2;84;57;50m-\033[38;2;82;56;49m_\033[38;2;81;57;49m_\033[38;2;81;58;50m-\033[38;2;82;60;51m-\033[38;2;84;63;53m-\033[38;2;87;66;56m?\033[38;2;91;71;57m1\033[38;2;96;76;59mt\033[38;2;94;76;57m1\033[38;2;106;94;81mr\033[38;2;202;200;198mh\033[38;2;255;255;255m$\033[0m                                                    \033[0m");
  $display("\033[0m                       \033[38;2;255;255;255m$\033[38;2;241;241;242m%%\033[38;2;158;155;153m0\033[38;2;91;80;71mt\033[38;2;79;62;47m_\033[38;2;76;54;42m+\033[38;2;86;62;51m-\033[38;2;87;64;52m-\033[38;2;86;62;50m-\033[38;2;86;60;50m-\033[38;2;85;60;51m-\033[38;2;82;58;49m-\033[38;2;86;57;48m-\033[38;2;80;53;47m_\033[38;2;80;54;49m_\033[38;2;109;68;60mt\033[38;2;117;76;67mj\033[38;2;147;93;83mu\033[38;2;136;93;83mu\033[38;2;97;64;55m1\033[38;2;103;70;60mt\033[38;2;105;83;75mj\033[38;2;135;117;108mz\033[38;2;144;126;117mY\033[38;2;151;136;126mJ\033[38;2;157;144;134mL\033[38;2;164;150;141mQ\033[38;2;172;158;148mO\033[38;2;168;154;144m0\033[38;2;156;141;132mC\033[38;2;118;102;94mu\033[38;2;96;68;58m1\033[38;2;100;69;58m1\033[38;2;90;63;55m?\033[38;2;99;65;57m1\033[38;2;90;58;49m-\033[38;2;85;57;49m-\033[38;2;84;57;50m-\033[38;2;77;55;48m_\033[38;2;71;52;47m+\033[38;2;82;57;50m-\033[38;2;80;57;49m_\033[38;2;78;58;49m_\033[38;2;79;59;51m-\033[38;2;82;61;52m-\033[38;2;85;62;54m-\033[38;2;86;65;55m?\033[38;2;87;68;54m?\033[38;2;85;70;54m?\033[38;2;96;86;75mf\033[38;2;141;138;135mJ\033[38;2;225;225;226mW\033[38;2;255;255;255m$$\033[0m                                                    \033[0m");
  $display("\033[0m                        \033[38;2;255;255;255m$$\033[38;2;215;215;217m*\033[38;2;156;152;148mQ\033[38;2;93;80;69mt\033[38;2;72;53;38m+\033[38;2;85;65;50m-\033[38;2;88;68;54m?\033[38;2;84;64;54m-\033[38;2;83;61;51m-\033[38;2;83;59;50m-\033[38;2;85;59;50m-\033[38;2;68;51;45m+\033[38;2;77;54;48m_\033[38;2;83;57;49m-\033[38;2;81;56;48m_\033[38;2;81;55;47m_\033[38;2;85;57;49m-\033[38;2;93;63;55m?\033[38;2;95;65;57m1\033[38;2;97;66;58m1\033[38;2;95;70;63m1\033[38;2;92;75;70mt\033[38;2;101;89;84mr\033[38;2;170;159;154mO\033[38;2;133;120;116mX\033[38;2;91;70;63m1\033[38;2;94;67;61m1\033[38;2;95;65;58m1\033[38;2;92;64;55m?\033[38;2;94;67;57m1\033[38;2;90;63;55m?\033[38;2;86;60;53m-\033[38;2;84;59;52m-\033[38;2;83;59;52m-\033[38;2;81;59;51m-\033[38;2;80;59;50m-\033[38;2;74;56;48m_\033[38;2;66;52;47m+\033[38;2;80;59;52m-\033[38;2;78;58;51m_\033[38;2;79;60;53m-\033[38;2;81;62;54m-\033[38;2;82;62;51m-\033[38;2;79;60;46m_\033[38;2;74;57;42m+\033[38;2;87;77;65m1\033[38;2;143;141;137mC\033[38;2;214;215;215m*\033[38;2;255;255;255m$$\033[0m                                                      \033[0m");
  $display("\033[0m                          \033[38;2;255;255;255m$$\033[38;2;222;223;223mM\033[38;2;142;138;134mJ\033[38;2;78;68;57m-\033[38;2;77;62;47m_\033[38;2;88;70;56m?\033[38;2;85;65;54m?\033[38;2;84;62;51m-\033[38;2;81;59;50m-\033[38;2;66;51;46m+\033[38;2;82;58;50m-\033[38;2;81;58;50m-\033[38;2;82;58;51m-\033[38;2;85;60;53m-\033[38;2;88;61;54m-\033[38;2;90;66;61m1\033[38;2;100;83;79mj\033[38;2;117;108;105mv\033[38;2;155;150;148mQ\033[38;2;208;206;205ma\033[38;2;172;169;168mm\033[38;2;245;242;240m%%\033[38;2;176;174;172mw\033[38;2;206;204;202ma\033[38;2;155;151;150mQ\033[38;2;135;127;125mY\033[38;2;112;96;92mn\033[38;2;94;73;65mt\033[38;2;88;65;56m?\033[38;2;84;62;55m-\033[38;2;82;61;54m-\033[38;2;80;60;53m-\033[38;2;78;60;52m-\033[38;2;77;60;52m-\033[38;2;74;58;50m_\033[38;2;64;52;46m+\033[38;2;80;62;52m-\033[38;2;79;61;52m-\033[38;2;76;58;49m_\033[38;2;70;53;40m+\033[38;2;67;51;35m~\033[38;2;86;75;63m1\033[38;2;150;147;142mL\033[38;2;213;214;214m*\033[38;2;255;255;255m$$\033[0m                                                        \033[0m");
  $display("\033[0m                            \033[38;2;255;255;255m$$\033[38;2;206;207;208mo\033[38;2;132;130;127mY\033[38;2;77;68;57m-\033[38;2;73;56;42m+\033[38;2;85;64;51m-\033[38;2;75;58;49m_\033[38;2;72;56;49m_\033[38;2;81;61;52m-\033[38;2;81;60;53m-\033[38;2;84;62;55m-\033[38;2;81;62;57m-\033[38;2;98;86;85mj\033[38;2;147;143;141mC\033[38;2;194;191;189mb\033[38;2;238;234;232m8\033[38;2;249;244;242mB\033[38;2;207;203;201ma\033[38;2;145;142;141mC\033[38;2;120;102;98mu\033[38;2;108;101;99mn\033[38;2;211;207;205mo\033[38;2;254;250;248m@\033[38;2;235;231;229m&\033[38;2;191;188;187md\033[38;2;163;159;157mO\033[38;2;125;117;114mz\033[38;2;89;74;69mt\033[38;2;82;61;54m-\033[38;2;79;61;54m-\033[38;2;76;61;52m-\033[38;2;77;60;52m-\033[38;2;76;61;52m-\033[38;2;62;53;47m+\033[38;2;69;55;46m+\033[38;2;62;48;37mi\033[38;2;59;47;34mi\033[38;2;88;79;68mt\033[38;2;158;154;150m0\033[38;2;220;222;222mM\033[38;2;255;255;255m$$\033[0m                                                          \033[0m");
  $display("\033[0m                              \033[38;2;255;255;255m$$\033[38;2;209;209;210mo\033[38;2;135;132;130mU\033[38;2;72;58;49m_\033[38;2;61;48;41m~\033[38;2;80;63;54m-\033[38;2;81;63;53m-\033[38;2;81;61;53m-\033[38;2;83;63;55m-\033[38;2;83;75;73mt\033[38;2;197;193;193mk\033[38;2;251;246;244mB\033[38;2;239;232;231m8\033[38;2;186;177;175mq\033[38;2;111;105;104mu\033[38;2;202;199;198mh\033[38;2;146;137;136mJ\033[38;2;103;73;65mt\033[38;2;140;130;126mU\033[38;2;219;216;215m#\033[38;2;143;138;136mJ\033[38;2;203;196;193mk\033[38;2;244;241;237m%%\033[38;2;252;249;245m@\033[38;2;220;218;217m#\033[38;2;107;101;100mn\033[38;2;78;58;52m_\033[38;2;80;62;54m-\033[38;2;76;61;53m-\033[38;2;78;60;51m-\033[38;2;78;63;53m-\033[38;2;72;60;52m_\033[38;2;55;46;39mi\033[38;2;84;78;70mt\033[38;2;163;161;158mO\033[38;2;227;227;227mW\033[38;2;255;255;255m$$\033[0m                                                            \033[0m");
  $display("\033[0m                                \033[38;2;255;255;255m$$\033[38;2;215;216;217m#\033[38;2;86;78;75mt\033[38;2;88;66;54m?\033[38;2;81;63;53m-\033[38;2;80;61;52m-\033[38;2;84;63;54m-\033[38;2;85;65;57m?\033[38;2;99;82;78mj\033[38;2;125;112;109mc\033[38;2;102;82;79mj\033[38;2;86;62;58m?\033[38;2;149;141;139mC\033[38;2;239;235;232m8\033[38;2;100;82;80mj\033[38;2;102;75;67mf\033[38;2;135;127;123mY\033[38;2;255;255;255m$\033[38;2;141;132;130mU\033[38;2;93;68;63m1\033[38;2;114;97;93mn\033[38;2;140;130;126mU\033[38;2;117;103;100mu\033[38;2;86;65;60m?\033[38;2;84;63;55m-\033[38;2;78;61;53m-\033[38;2;77;61;52m-\033[38;2;79;62;52m-\033[38;2;82;64;54m-\033[38;2;87;68;56m?\033[38;2;116;111;107mv\033[38;2;236;237;237m8\033[38;2;255;255;255m$$\033[0m                                                              \033[0m");
  $display("\033[0m                                 \033[38;2;255;255;255m$\033[38;2;240;241;241m%%\033[38;2;102;88;79mj\033[38;2;92;68;55m?\033[38;2;83;63;53m-\033[38;2;80;60;53m-\033[38;2;79;60;52m-\033[38;2;80;60;53m-\033[38;2;82;59;53m-\033[38;2;83;58;52m-\033[38;2;94;67;61m1\033[38;2;88;74;71mt\033[38;2;236;229;227m&\033[38;2;169;161;160mZ\033[38;2;92;67;62m1\033[38;2;102;71;66mt\033[38;2;109;96;94mn\033[38;2;253;248;246m@\033[38;2;180;174;173mw\033[38;2;85;64;62m?\033[38;2;92;67;62m1\033[38;2;81;58;53m-\033[38;2;79;59;53m-\033[38;2;81;62;56m-\033[38;2;79;61;54m-\033[38;2;77;61;53m--\033[38;2;79;62;52m-\033[38;2;83;65;54m-\033[38;2;93;72;59m1\033[38;2;123;114;107mc\033[38;2;252;253;255m$\033[38;2;255;255;255m$\033[0m                                                               \033[0m");
  $display("\033[0m                                 \033[38;2;255;255;255m$\033[38;2;206;205;203ma\033[38;2;97;74;59m1\033[38;2;93;68;57m1\033[38;2;83;62;53m-\033[38;2;80;60;51m-\033[38;2;78;60;51m-\033[38;2;78;59;51m_\033[38;2;79;60;54m-\033[38;2;86;64;58m?\033[38;2;83;61;56m-\033[38;2;133;128;126mY\033[38;2;249;242;241mB\033[38;2;101;87;85mr\033[38;2;99;69;63mt\033[38;2;99;71;65mt\033[38;2;90;73;70mt\033[38;2;223;218;215m#\033[38;2;231;226;224mW\033[38;2;87;73;73mt\033[38;2;88;67;62m1\033[38;2;82;63;57m-\033[38;2;78;60;54m-\033[38;2;77;59;55m-\033[38;2;76;61;54m-\033[38;2;76;61;52m-\033[38;2;75;61;50m_\033[38;2;77;61;51m-\033[38;2;82;64;53m-\033[38;2;96;75;61mt\033[38;2;89;74;61m1\033[38;2;209;210;210mo\033[38;2;255;255;255m$\033[0m                                                               \033[0m");
  $display("\033[0m                                \033[38;2;255;255;255m$$\033[38;2;139;133;126mU\033[38;2;97;72;56m1\033[38;2;89;67;56m?\033[38;2;81;61;50m-\033[38;2;79;60;49m_\033[38;2;78;59;52m-\033[38;2;77;60;53m-\033[38;2;79;61;55m-\033[38;2;88;65;58m?\033[38;2;85;72;68m1\033[38;2;226;221;219mM\033[38;2;199;194;192mk\033[38;2;81;61;57m-\033[38;2;95;68;62m1\033[38;2;93;68;63m1\033[38;2;82;63;59m?\033[38;2;178;172;171mw\033[38;2;255;253;252m$\033[38;2;122;112;112mc\033[38;2;87;62;60m?\033[38;2;84;63;58m?\033[38;2;77;59;56m-\033[38;2;76;59;55m-\033[38;2;77;60;52m-\033[38;2;78;60;51m-\033[38;2;77;61;51m--\033[38;2;81;64;53m-\033[38;2;92;71;59m1\033[38;2;92;71;57m1\033[38;2;138;137;136mJ\033[38;2;255;255;255m$\033[0m                                                               \033[0m");
  $display("\033[0m                                \033[38;2;255;255;255m$\033[38;2;242;243;243m%%\033[38;2;115;101;87mn\033[38;2;96;72;57m1\033[38;2;85;65;54m?\033[38;2;80;60;50m-\033[38;2;79;60;50m-\033[38;2;76;60;52m_\033[38;2;76;60;53m-\033[38;2;80;62;56m-\033[38;2;78;58;53m-\033[38;2;140;134;132mJ\033[38;2;255;255;255m$\033[38;2;154;147;146mQ\033[38;2;81;56;50m_\033[38;2;86;64;58m?\033[38;2;86;65;59m?\033[38;2;84;62;57m-\033[38;2;136;129;127mY\033[38;2;255;255;254m$\033[38;2;182;176;173mq\033[38;2;80;58;56m-\033[38;2;85;64;58m?\033[38;2;78;60;55m-\033[38;2;76;59;53m_\033[38;2;76;59;51m__\033[38;2;77;61;51m-\033[38;2;78;61;51m-\033[38;2;80;62;51m-\033[38;2;88;68;56m?\033[38;2;99;75;60mt\033[38;2;111;105;99mu\033[38;2;251;252;252m@\033[38;2;255;255;255m$\033[0m                                                              \033[0m");
  $display("\033[0m                                \033[38;2;255;255;255m$\033[38;2;219;218;216m#\033[38;2;110;87;67mj\033[38;2;93;69;55m1\033[38;2;83;63;54m-\033[38;2;79;61;51m-\033[38;2;77;59;51m_\033[38;2;75;58;51m_\033[38;2;74;59;53m_\033[38;2;78;61;56m-\033[38;2;75;57;51m_\033[38;2;138;130;128mU\033[38;2;211;207;206mo\033[38;2;102;91;88mr\033[38;2;84;58;55m-\033[38;2;81;60;56m-\033[38;2;80;62;56m-\033[38;2;86;63;60m?\033[38;2;86;72;71m1\033[38;2;228;222;217mM\033[38;2;229;223;218mM\033[38;2;89;76;74mt\033[38;2;83;61;55m-\033[38;2;78;60;55m-\033[38;2;76;58;52m_\033[38;2;76;58;51m_\033[38;2;76;59;51m_\033[38;2;76;60;51m_\033[38;2;78;61;51m-\033[38;2;79;61;51m-\033[38;2;86;66;53m?\033[38;2;101;78;62mt\033[38;2;88;78;67mt\033[38;2;222;223;224mM\033[38;2;255;255;255m$\033[0m                                                              \033[0m");
  $display("\033[0m                               \033[38;2;255;255;255m$$\033[38;2;150;142;135mC\033[38;2;96;67;49m?\033[38;2;85;60;49m-\033[38;2;76;55;46m_\033[38;2;71;54;44m+\033[38;2;70;53;44m+\033[38;2;68;52;43m+\033[38;2;66;52;43m~\033[38;2;69;52;45m+\033[38;2;74;54;47m+\033[38;2;70;52;44m+\033[38;2;70;52;46m+\033[38;2;72;52;46m+\033[38;2;74;53;48m+\033[38;2;72;52;48m+\033[38;2;72;53;48m+\033[38;2;74;54;50m_\033[38;2;74;54;51m_\033[38;2;92;78;75mf\033[38;2;93;77;74mf\033[38;2;75;56;53m_\033[38;2;73;53;48m+\033[38;2;72;53;46m+\033[38;2;71;53;45m+++\033[38;2;72;54;46m+\033[38;2;73;55;46m+\033[38;2;75;55;46m+\033[38;2;78;58;46m_\033[38;2;91;70;54m?\033[38;2;79;64;47m-\033[38;2;168;168;168mm\033[38;2;255;255;255m$\033[0m                                                              \033[0m");
  $display("\033[0m                               \033[38;2;255;255;255m$\033[38;2;253;253;253m$\033[38;2;194;184;176mp\033[38;2;172;156;149mO\033[38;2;166;153;148m0\033[38;2;163;151;147m0\033[38;2;159;151;146mQ\033[38;2;158;150;146mQQ\033[38;2;157;150;146mQQ\033[38;2;158;149;146mQ\033[38;2;159;149;147mQ\033[38;2;159;149;146mQ\033[38;2;159;149;147mQQ\033[38;2;159;150;148mQQQ\033[38;2;160;151;148m0\033[38;2;158;148;146mQQ\033[38;2;160;151;148m0\033[38;2;159;150;148mQ\033[38;2;159;151;147mQQQQ\033[38;2;160;151;147mQQ\033[38;2;161;152;147m0\033[38;2;163;153;148m0\033[38;2;167;157;151mO\033[38;2;171;160;150mO\033[38;2;201;199;197mh\033[38;2;255;255;255m$\033[0m                                                              \033[0m");
  $display("\033[0m                                \033[38;2;255;255;255m$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$\033[0m                                                              \033[0m");
  $display ("--------------------------------------------------");
  $display("                  Congratulations!               ");
  $display("              execution cycles = %7d", total_latency);
  $display("              clock period = %4fns", CYCLE);
  $display ("--------------------------------------------------");
  $finish;	
endtask

task fail_task;
  $display("\033[0m                                                \033[38;2;255;255;255m$$$\033[38;2;247;247;247mB\033[38;2;241;241;241m%%\033[38;2;252;252;252m$\033[38;2;255;255;255m$$$\033[0m                                          \033[0m");
  $display("\033[0m                                             \033[38;2;255;255;255m$$\033[38;2;226;226;228mW\033[38;2;162;163;170mZ\033[38;2;116;119;128mz\033[38;2;98;102;113mu\033[38;2;95;99;112mn\033[38;2;94;98;111mn\033[38;2;93;96;107mx\033[38;2;95;99;106mn\033[38;2;122;125;127mX\033[38;2;167;167;169mm\033[38;2;231;231;229m&\033[38;2;255;255;255m$\033[0m                                        \033[0m");
  $display("\033[0m                                            \033[38;2;255;255;255m$\033[38;2;223;229;229mW\033[38;2;132;138;145mJ\033[38;2;60;66;81m?\033[38;2;72;77;91mt\033[38;2;107;112;123mc\033[38;2;145;148;157mQ\033[38;2;173;175;181mq\033[38;2;188;190;196mb\033[38;2;186;187;193md\033[38;2;123;126;137mY\033[38;2;30;36;53ml\033[38;2;30;35;52ml\033[38;2;67;71;85m1\033[38;2;159;158;161mO\033[38;2;251;251;248m@\033[38;2;255;255;255m$\033[0m                                      \033[0m");
  $display("\033[0m                                          \033[38;2;255;0;0mf\033[38;2;255;59;59mX\033[38;2;234;163;162md\033[38;2;110;60;68mt\033[38;2;80;57;69m?\033[38;2;189;197;202mk\033[38;2;249;255;253m$\033[38;2;255;255;255m$$$$$$\033[38;2;186;187;192md\033[38;2;37;43;58mi\033[38;2;30;36;54ml\033[38;2;27;30;45mI\033[38;2;189;186;184md\033[38;2;255;255;255m$\033[0m                                      \033[0m");
  $display("\033[0m                                \033[38;2;255;0;0mfffffff\033[38;2;255;1;1mf\033[38;2;255;2;2mj\033[38;2;255;0;0mff\033[38;2;255;69;69mU\033[38;2;254;65;65mY\033[38;2;249;51;52mz\033[38;2;255;34;33mu\033[38;2;244;84;86mJ\033[38;2;126;111;134mX\033[38;2;100;118;147mz\033[38;2;107;123;150mY\033[38;2;104;119;147mX\033[38;2;106;120;146mX\033[38;2;95;109;130mv\033[38;2;90;100;112mn\033[38;2;111;114;121mc\033[38;2;39;45;57mi\033[38;2;33;39;56m!\033[38;2;28;33;50ml\033[38;2;122;126;131mY\033[38;2;179;187;188mp\033[38;2;192;195;195mk\033[38;2;224;224;224mM\033[38;2;255;255;252m$\033[38;2;255;255;255m$\033[0m                                  \033[0m");
  $display("\033[0m                     \033[38;2;255;0;0mffff\033[0m    \033[38;2;255;0;0mfff\033[38;2;255;11;11mr\033[38;2;255;38;38mv\033[38;2;255;79;79mJ\033[38;2;255;109;109m0\033[38;2;255;141;141mq\033[38;2;255;173;173mh\033[38;2;255;195;195m*\033[38;2;255;210;210mW\033[38;2;255;215;215mW\033[38;2;255;154;154md\033[38;2;255;57;57mX\033[38;2;255;235;235m%%\033[38;2;255;255;255m$$\033[38;2;255;180;180ma\033[38;2;255;0;0mf\033[38;2;169;29;46mf\033[38;2;46;80;121mf\033[38;2;52;75;111mt\033[38;2;50;74;108mt\033[38;2;50;73;106m1\033[38;2;47;71;104m1\033[38;2;40;62;91m-\033[38;2;28;45;69mi\033[38;2;28;38;58m!\033[38;2;30;36;53ml\033[38;2;32;39;57m!\033[38;2;30;42;60m!\033[38;2;32;47;63mi\033[38;2;44;60;77m_\033[38;2;68;83;100mf\033[38;2;105;115;128mc\033[38;2;154;160;162mO\033[38;2;211;211;211mo\033[38;2;255;255;255m$$\033[0m                               \033[0m");
  $display("\033[0m           \033[38;2;255;0;0mffffff\033[0m   \033[38;2;255;0;0mff\033[38;2;255;21;21mn\033[38;2;255;14;14mr\033[38;2;255;2;2mj\033[38;2;255;0;0mff\033[0m  \033[38;2;255;0;0mff\033[38;2;255;143;143mp\033[38;2;255;225;225m8\033[38;2;255;252;252m$\033[38;2;255;255;255m$$$$\033[38;2;255;248;248m@\033[38;2;255;223;223m&\033[38;2;255;189;188mo\033[38;2;255;138;138mq\033[38;2;255;100;100mQ\033[38;2;255;251;251m$\033[38;2;255;255;255m$$\033[38;2;255;154;154md\033[38;2;255;0;0mf\033[38;2;127;49;72mf\033[38;2;48;81;119mf\033[38;2;54;80;115mf\033[38;2;50;79;113mt\033[38;2;51;75;108mt\033[38;2;53;73;107mt\033[38;2;54;74;109mt\033[38;2;52;74;109mt\033[38;2;47;67;101m?\033[38;2;35;49;71m~\033[38;2;27;36;51ml\033[38;2;27;36;50ml\033[38;2;28;36;52ml\033[38;2;26;35;53ml\033[38;2;25;34;53ml\033[38;2;25;34;54ml\033[38;2;29;44;62mi\033[38;2;56;72;87m?\033[38;2;116;127;136mY\033[38;2;190;192;194mb\033[38;2;255;255;255m$$\033[0m                             \033[0m");
  $display("\033[0m       \033[38;2;255;0;0mffff\033[38;2;255;15;15mx\033[38;2;255;45;45mc\033[38;2;255;77;77mJ\033[38;2;255;101;101mQ\033[38;2;255;79;79mJ\033[38;2;255;22;22mn\033[38;2;255;0;0mffff\033[38;2;255;110;110mO\033[38;2;255;233;233m%%\033[38;2;255;224;224m8\033[38;2;255;202;202m#\033[38;2;255;43;43mc\033[38;2;255;0;0mff\033[0m \033[38;2;255;0;0mff\033[38;2;255;70;70mU\033[38;2;255;210;210mWW\033[38;2;255;158;158mb\033[38;2;255;236;236m%%\033[38;2;255;255;255m$$\033[38;2;255;79;79mJ\033[38;2;248;9;10mj\033[38;2;225;9;15mf\033[38;2;255;0;0mf\033[38;2;255;131;131mw\033[38;2;255;255;255m$$\033[38;2;255;254;254m$\033[38;2;255;67;67mY\033[38;2;240;1;3mf\033[38;2;74;76;109mj\033[38;2;53;81;118mf\033[38;2;51;77;111mt\033[38;2;52;77;110mt\033[38;2;55;78;111mf\033[38;2;56;79;111mf\033[38;2;55;79;111mf\033[38;2;54;78;111mf\033[38;2;53;77;112mt\033[38;2;54;76;111mt\033[38;2;44;62;88m-\033[38;2;29;42;58m!\033[38;2;27;36;52ml\033[38;2;29;37;53ml\033[38;2;28;36;54ml\033[38;2;28;36;53ml\033[38;2;27;33;51ml\033[38;2;24;34;51ml\033[38;2;27;42;61m!\033[38;2;46;61;80m_\033[38;2;114;121;129mz\033[38;2;202;201;202mh\033[38;2;255;255;255m$$\033[0m                           \033[0m");
  $display("\033[0m    \033[38;2;255;0;0mfff\033[38;2;255;8;8mr\033[38;2;255;51;51mz\033[38;2;255;113;113mO\033[38;2;255;178;178ma\033[38;2;255;228;228m8\033[38;2;255;255;255m$$$$\033[38;2;255;222;222m&\033[38;2;255;58;58mX\033[38;2;255;4;4mj\033[38;2;255;84;84mC\033[38;2;255;153;153md\033[38;2;255;253;253m$\033[38;2;255;255;255m$$$\033[38;2;255;186;186mo\033[38;2;255;3;3mj\033[38;2;255;0;0mf\033[0m  \033[38;2;255;0;0mf\033[38;2;255;37;37mv\033[38;2;252;48;47mc\033[38;2;250;6;7mj\033[38;2;255;12;12mr\033[38;2;255;233;233m%%\033[38;2;255;255;255m$\033[38;2;255;246;246m@\033[38;2;255;31;30mu\033[38;2;208;14;23mf\033[38;2;169;37;54mj\033[38;2;255;2;2mj\033[38;2;255;203;203m#\033[38;2;255;255;255m$$\033[38;2;255;226;226m8\033[38;2;255;10;9mr\033[38;2;186;25;37mf\033[38;2;38;83;118mt\033[38;2;46;78;111mt\033[38;2;54;77;110mt\033[38;2;58;77;111mf\033[38;2;53;80;114mf\033[38;2;47;81;118mff\033[38;2;51;78;112mt\033[38;2;54;77;111mt\033[38;2;53;76;113mt\033[38;2;53;75;111mt\033[38;2;48;70;100m1\033[38;2;31;45;68mi\033[38;2;26;33;49ml\033[38;2;25;35;52ml\033[38;2;27;33;52ml\033[38;2;28;31;50ml\033[38;2;28;31;51ml\033[38;2;27;31;50ml\033[38;2;28;38;55ml\033[38;2;33;50;66mi\033[38;2;53;70;85m?\033[38;2;142;146;149mL\033[38;2;234;234;232m&\033[38;2;255;255;255m$\033[0m                          \033[0m");
  $display("\033[0m  \033[38;2;255;0;0mff\033[38;2;255;22;22mn\033[38;2;255;75;75mJ\033[38;2;255;149;149mp\033[38;2;255;214;214mW\033[38;2;255;253;253m$\033[38;2;255;255;255m$$\033[38;2;255;236;236m%%\033[38;2;255;191;191m*\033[38;2;255;143;143mp\033[38;2;255;100;100mQ\033[38;2;255;68;68mY\033[38;2;255;46;46mc\033[38;2;255;7;7mj\033[38;2;255;115;115mO\033[38;2;255;255;255m$$$\033[38;2;255;249;249m@\033[38;2;255;255;255m$$$\033[38;2;255;117;117mZ\033[38;2;255;0;0mfff\033[38;2;255;214;214mW\033[38;2;202;218;222m*\033[38;2;119;115;134mX\033[38;2;231;1;5mt\033[38;2;255;53;53mz\033[38;2;255;254;254m$\033[38;2;255;255;255m$\033[38;2;255;220;220m&\033[38;2;255;6;5mj\033[38;2;184;29;43mf\033[38;2;214;13;21mf\033[38;2;255;37;36mv\033[38;2;255;247;247m@\033[38;2;255;255;255m$$\033[38;2;255;156;156mb\033[38;2;255;0;0mf\033[38;2;193;11;21m1\033[38;2;161;25;40m1\033[38;2;192;20;31mf\033[38;2;213;19;27mj\033[38;2;216;19;26mj\033[38;2;196;17;28mt\033[38;2;166;24;42mt\033[38;2;134;42;67mf\033[38;2;71;69;104mf\033[38;2;49;77;114mt\033[38;2;52;74;109mt\033[38;2;51;74;108mtt\033[38;2;50;72;105m1\033[38;2;34;47;70m~\033[38;2;27;32;51ml\033[38;2;26;35;53ml\033[38;2;25;36;52ml\033[38;2;27;34;52ml\033[38;2;26;32;50ml\033[38;2;26;30;49mI\033[38;2;25;32;48mI\033[38;2;33;50;64mi\033[38;2;36;57;73m+\033[38;2;84;95;106mx\033[38;2;202;204;203ma\033[38;2;255;255;255m$\033[0m                         \033[0m");
  $display("\033[0m  \033[38;2;255;0;0mf\033[38;2;255;6;6mj\033[38;2;255;195;195m*\033[38;2;255;255;255m$$$$\033[38;2;255;212;212mW\033[38;2;255;71;71mU\033[38;2;255;18;18mx\033[38;2;255;0;0mfffff\033[38;2;255;21;21mn\033[38;2;255;232;232m%%\033[38;2;255;255;255m$$\033[38;2;255;238;238mB\033[38;2;255;62;62mY\033[38;2;255;130;130mw\033[38;2;255;253;253m$\033[38;2;255;255;255m$\033[38;2;255;247;247m@\033[38;2;255;121;121mZ\033[38;2;255;103;103m0\033[38;2;255;65;65mY\033[38;2;255;35;35mv\033[38;2;187;38;49mr\033[38;2;116;55;81mf\033[38;2;255;0;0mf\033[38;2;255;137;137mq\033[38;2;255;255;255m$$\033[38;2;255;181;181ma\033[38;2;255;0;0mf\033[38;2;179;29;44mf\033[38;2;234;1;5mt\033[38;2;255;78;78mJ\033[38;2;255;255;255m$$$\033[38;2;255;121;121mZ\033[38;2;255;47;47mc\033[38;2;255;105;104m0\033[38;2;255;147;145mp\033[38;2;255;179;178ma\033[38;2;255;206;205mM\033[38;2;255;211;210mW\033[38;2;255;180;179ma\033[38;2;255;149;148mp\033[38;2;255;35;33mu\033[38;2;215;14;22mf\033[38;2;67;68;101mt\033[38;2;45;71;104m1\033[38;2;53;75;110mt\033[38;2;52;75;108mt\033[38;2;51;75;107mt\033[38;2;50;71;103m1\033[38;2;34;46;70m~\033[38;2;25;34;51ml\033[38;2;25;37;54ml\033[38;2;25;35;52mll\033[38;2;25;33;50ml\033[38;2;25;32;49mI\033[38;2;23;30;48mI\033[38;2;35;46;63mi\033[38;2;38;59;76m+\033[38;2;55;73;87m?\033[38;2;177;182;184mp\033[38;2;255;255;255m$\033[0m                        \033[0m");
  $display("\033[0m  \033[38;2;255;0;0mff\033[38;2;255;43;43mc\033[38;2;255;141;141mq\033[38;2;255;233;233m%%\033[38;2;255;255;255m$$\033[38;2;255;127;127mm\033[38;2;255;0;0mf\033[38;2;255;5;5mj\033[38;2;255;33;33mu\033[38;2;255;58;58mX\033[38;2;255;26;26mn\033[38;2;255;1;1mf\033[38;2;255;0;0mf\033[38;2;255;106;106m0\033[38;2;255;255;255m$$$\033[38;2;255;139;139mq\033[38;2;255;58;58mX\033[38;2;255;114;114mO\033[38;2;255;245;245m@\033[38;2;255;255;255m$$$$\033[38;2;255;188;188mo\033[38;2;255;15;14mr\033[38;2;229;1;6mt\033[38;2;206;11;20mt\033[38;2;255;6;5mj\033[38;2;255;219;219m&\033[38;2;255;255;255m$$\033[38;2;255;137;137mq\033[38;2;255;51;51mz\033[38;2;246;22;23mx\033[38;2;253;1;1mf\033[38;2;255;54;54mz\033[38;2;255;254;254m$\033[38;2;255;255;255m$$\033[38;2;255;248;248m@\033[38;2;255;254;254m$\033[38;2;255;255;255m$$$$\033[38;2;255;245;245m@\033[38;2;255;242;242mB\033[38;2;255;223;223m&\033[38;2;255;90;89mL\033[38;2;255;0;0mf\033[38;2;112;46;69m1\033[38;2;43;75;109m1\033[38;2;54;77;111mt\033[38;2;53;76;110mt\033[38;2;52;75;108mt\033[38;2;51;74;108mt\033[38;2;49;70;103m1\033[38;2;28;41;62m!\033[38;2;26;33;51ml\033[38;2;26;34;53ml\033[38;2;26;35;52mll\033[38;2;26;34;51ml\033[38;2;26;32;51ml\033[38;2;25;28;43mI\033[38;2;35;45;62mi\033[38;2;39;62;80m_\033[38;2;46;64;81m-\033[38;2;171;176;178mw\033[38;2;255;255;255m$\033[0m                       \033[0m");
  $display("\033[0m \033[38;2;255;0;0mff\033[38;2;255;1;1mf\033[38;2;255;37;37mv\033[38;2;255;54;54mz\033[38;2;255;219;219m&\033[38;2;255;255;255m$$\033[38;2;255;190;190mo\033[38;2;255;178;178ma\033[38;2;255;222;222m&\033[38;2;255;251;251m$\033[38;2;255;255;255m$\033[38;2;255;213;213mW\033[38;2;255;19;19mx\033[38;2;255;10;10mr\033[38;2;255;218;218m&\033[38;2;255;255;255m$$\033[38;2;255;250;250m@\033[38;2;255;252;252m$\033[38;2;255;255;255m$$$\033[38;2;255;240;240mB\033[38;2;255;255;255m$$\033[38;2;255;238;238mB\033[38;2;255;35;35mv\033[38;2;255;17;17mx\033[38;2;254;53;54mz\033[38;2;255;95;94mL\033[38;2;255;162;162mb\033[38;2;255;255;255m$$$$$\033[38;2;255;227;226m8\033[38;2;255;52;52mz\033[38;2;255;0;0mf\033[38;2;255;96;95mL\033[38;2;255;229;229m8\033[38;2;255;255;255m$$\033[38;2;255;240;239mB\033[38;2;255;195;194m*\033[38;2;255;130;129mw\033[38;2;255;83;83mC\033[38;2;251;49;49mc\033[38;2;237;32;33mn\033[38;2;234;30;33mn\033[38;2;223;20;25mj\033[38;2;192;20;31mf\033[38;2;120;46;68mt\033[38;2;81;82;95mj\033[38;2;54;75;105mt\033[38;2;54;76;112mt\033[38;2;53;77;112mt\033[38;2;53;75;110mt\033[38;2;52;74;106mt\033[38;2;53;75;108mt\033[38;2;44;63;88m-\033[38;2;24;36;53ml\033[38;2;27;37;53ml\033[38;2;26;35;52ml\033[38;2;25;34;51ml\033[38;2;26;35;52ml\033[38;2;25;34;51ml\033[38;2;25;32;49mI\033[38;2;25;30;46mI\033[38;2;36;49;66m~\033[38;2;40;63;80m_\033[38;2;44;63;78m_\033[38;2;171;175;177mw\033[38;2;255;255;255m$\033[0m                      \033[0m");
  $display("\033[0m \033[38;2;255;0;0mff\033[38;2;255;89;89mL\033[38;2;255;255;255m$$$$$$$\033[38;2;255;227;227m8\033[38;2;255;187;187mo\033[38;2;255;135;135mw\033[38;2;255;66;66mY\033[38;2;255;0;0mf\033[38;2;255;99;99mQ\033[38;2;255;255;255m$$\033[38;2;255;247;247m@\033[38;2;255;84;84mC\033[38;2;255;141;141mq\033[38;2;255;161;161mb\033[38;2;255;118;118mZ\033[38;2;255;77;77mJ\033[38;2;255;132;132mw\033[38;2;255;255;255m$$$\033[38;2;255;70;70mU\033[38;2;255;110;110mO\033[38;2;255;255;255m$$$\033[38;2;255;239;239mB\033[38;2;255;207;206mM\033[38;2;255;184;183mo\033[38;2;255;146;145mp\033[38;2;255;104;103m0\033[38;2;255;67;67mY\033[38;2;242;12;15mj\033[38;2;171;34;50mf\033[38;2;204;12;21mt\033[38;2;246;29;30mn\033[38;2;254;60;61mX\033[38;2;253;56;57mX\033[38;2;243;32;35mn\033[38;2;217;15;22mf\033[38;2;169;22;36m1\033[38;2;103;22;37m+\033[38;2;71;28;45mi\033[38;2;66;61;88m?\033[38;2;65;70;101mt\033[38;2;55;70;106mt\033[38;2;43;72;104m1\033[38;2;102;106;104mu\033[38;2;162;139;110mJ\033[38;2;61;77;97mt\033[38;2;53;73;103m1\033[38;2;55;73;102m1\033[38;2;52;76;111mt\033[38;2;52;75;108mt\033[38;2;49;72;104m1\033[38;2;47;68;101m1\033[38;2;34;46;69mi\033[38;2;26;36;52ml\033[38;2;27;37;54ml\033[38;2;24;31;49mI\033[38;2;25;33;51ml\033[38;2;25;34;51ml\033[38;2;25;35;52ml\033[38;2;26;32;50ml\033[38;2;25;32;47mI\033[38;2;37;54;69m~\033[38;2;39;61;77m_\033[38;2;45;64;80m-\033[38;2;200;202;202mh\033[38;2;255;255;255m$\033[0m                     \033[0m");
  $display("\033[0m \033[38;2;255;0;0mff\033[38;2;255;28;28mn\033[38;2;255;158;158mb\033[38;2;255;245;245m@\033[38;2;255;255;255m$$\033[38;2;255;189;189mo\033[38;2;255;90;90mL\033[38;2;255;43;43mc\033[38;2;255;13;13mr\033[38;2;255;0;0mfff\033[38;2;255;2;2mj\033[38;2;255;198;198m#\033[38;2;255;255;255m$$\033[38;2;255;204;204mM\033[38;2;255;0;0mfff\033[38;2;255;16;14mx\033[38;2;255;13;12mr\033[38;2;255;139;138mq\033[38;2;255;235;235m%%\033[38;2;255;224;223m8\033[38;2;255;124;122mm\033[38;2;255;4;4mj\033[38;2;255;8;8mr\033[38;2;255;112;111mO\033[38;2;255;126;125mm\033[38;2;255;74;73mU\033[38;2;246;33;35mu\033[38;2;218;19;26mj\033[38;2;193;21;33mf\033[38;2;185;20;34mt\033[38;2;138;38;59mt\033[38;2;111;52;79mt\033[38;2;83;70;103mf\033[38;2;49;82;121mf\033[38;2;49;70;107m1\033[38;2;74;57;88m1\033[38;2;92;52;79m1\033[38;2;91;58;85mt\033[38;2;76;65;98mt\033[38;2;57;76;111mf\033[38;2;34;61;87m_\033[38;2;22;41;61m!\033[38;2;45;69;97m?\033[38;2;50;77;113mt\033[38;2;44;71;109m1\033[38;2;61;75;97mt\033[38;2;133;123;102mz\033[38;2;207;181;139mw\033[38;2;220;193;156mb\033[38;2;88;89;98mr\033[38;2;55;74;94m1\033[38;2;115;108;101mv\033[38;2;51;71;98m1\033[38;2;52;74;107mt\033[38;2;53;73;104m1\033[38;2;37;54;83m+\033[38;2;40;56;82m_\033[38;2;27;35;52ml\033[38;2;25;37;54ml\033[38;2;25;33;49mI\033[38;2;23;32;47mI\033[38;2;26;34;52ml\033[38;2;26;34;51ml\033[38;2;26;33;51ml\033[38;2;25;30;47mI\033[38;2;26;36;52ml\033[38;2;37;60;74m+\033[38;2;34;55;76m+\033[38;2;80;92;102mr\033[38;2;237;237;234m8\033[38;2;255;255;255m$\033[0m                    \033[0m");
  $display("\033[0m  \033[38;2;255;0;0mfff\033[38;2;255;219;219m&\033[38;2;255;255;255m$$\033[38;2;255;69;69mU\033[38;2;255;0;0mfff\033[0m  \033[38;2;255;0;0mf\033[38;2;255;1;1mf\033[38;2;255;89;89mL\033[38;2;255;206;206mM\033[38;2;255;208;208mM\033[38;2;255;84;84mC\033[38;2;253;0;0mf\033[38;2;255;85;85mC\033[38;2;255;255;255m$\033[38;2;168;164;176mm\033[38;2;162;40;57mj\033[38;2;217;13;20mf\033[38;2;239;31;34mn\033[38;2;235;25;29mx\033[38;2;199;17;28mf\033[38;2;121;57;84mj\033[38;2;107;61;91mj\033[38;2;156;29;46mt\033[38;2;154;32;51mt\033[38;2;119;49;75mf\033[38;2;80;68;103mf\033[38;2;57;80;119mf\033[38;2;49;84;125mj\033[38;2;49;85;125mj\033[38;2;48;85;122mf\033[38;2;52;83;122mf\033[38;2;54;81;120mf\033[38;2;55;77;114mf\033[38;2;47;70;106m1\033[38;2;40;65;94m-\033[38;2;47;77;108mt\033[38;2;50;80;114mf\033[38;2;50;79;114mf\033[38;2;48;72;102m1\033[38;2;29;39;63m!\033[38;2;46;62;90m-\033[38;2;49;73;108m1\033[38;2;52;67;100m1\033[38;2;103;99;101mn\033[38;2;189;165;131mO\033[38;2;233;212;169ma\033[38;2;246;226;187m#\033[38;2;250;230;191mM\033[38;2;181;169;153mm\033[38;2;50;63;90m-\033[38;2;143;126;112mY\033[38;2;121;115;115mz\033[38;2;49;67;96m?\033[38;2;57;75;106mt\033[38;2;40;55;81m+\033[38;2;34;48;70m~\033[38;2;28;39;60m!\033[38;2;25;36;53ml\033[38;2;26;34;52ml\033[38;2;23;30;49mI\033[38;2;26;34;52ml\033[38;2;26;34;51ml\033[38;2;26;34;52ml\033[38;2;26;33;49ml\033[38;2;23;30;46mI\033[38;2;30;45;60mi\033[38;2;38;60;76m+\033[38;2;32;53;73m~\033[38;2;129;136;142mJ\033[38;2;255;255;255m$\033[0m                    \033[0m");
  $display("\033[0m   \033[38;2;255;0;0mf\033[38;2;255;1;1mf\033[38;2;255;113;113mO\033[38;2;255;227;227m8\033[38;2;255;237;237mB\033[38;2;255;63;63mY\033[38;2;255;0;0mff\033[0m    \033[38;2;255;0;0mff\033[38;2;255;4;4mj\033[38;2;255;2;2mj\033[38;2;255;0;0mf\033[38;2;255;163;160mb\033[38;2;216;225;229mM\033[38;2;117;132;156mJ\033[38;2;51;77;116mf\033[38;2;52;88;126mj\033[38;2;61;83;121mj\033[38;2;78;77;112mj\033[38;2;74;78;114mj\033[38;2;57;86;127mr\033[38;2;52;87;128mj\033[38;2;48;81;120mf\033[38;2;47;84;120mf\033[38;2;48;86;126mj\033[38;2;48;85;126mj\033[38;2;52;84;124mj\033[38;2;55;82;122mj\033[38;2;55;82;121mj\033[38;2;57;81;120mj\033[38;2;58;79;117mf\033[38;2;56;78;117mff\033[38;2;55;76;114mf\033[38;2;45;67;100m?\033[38;2;46;65;95m?\033[38;2;54;76;111mt\033[38;2;54;78;111mf\033[38;2;57;80;112mf\033[38;2;39;54;77m+\033[38;2;28;45;72mi\033[38;2;58;75;104mt\033[38;2;102;107;117mv\033[38;2;182;167;148mZ\033[38;2;237;217;179mo\033[38;2;246;231;195mM\033[38;2;248;230;195mM\033[38;2;247;228;192mM\033[38;2;248;229;193mM\033[38;2;251;232;199mW\033[38;2;125;126;128mY\033[38;2;94;88;90mr\033[38;2;210;188;155mp\033[38;2;83;90;105mr\033[38;2;49;69;101m1\033[38;2;46;64;90m-\033[38;2;29;39;59m!\033[38;2;30;40;58m!\033[38;2;27;37;55ml\033[38;2;28;37;55ml\033[38;2;25;30;50mI\033[38;2;25;33;50ml\033[38;2;27;36;53ml\033[38;2;26;35;52mll\033[38;2;24;32;49mI\033[38;2;24;33;51ml\033[38;2;37;55;73m+\033[38;2;39;59;78m+\033[38;2;39;56;73m+\033[38;2;177;180;182mq\033[38;2;255;255;255m$\033[0m                   \033[0m");
  $display("\033[0m    \033[38;2;255;0;0mff\033[38;2;255;19;19mx\033[38;2;255;27;27mn\033[38;2;255;0;0mfff\033[0m      \033[38;2;255;0;0mf\033[38;2;255;223;207mW\033[38;2;255;255;255m$\033[38;2;168;183;196mp\033[38;2;69;94;129mx\033[38;2;105;125;154mY\033[38;2;180;190;204mb\033[38;2;88;110;143mc\033[38;2;56;82;124mj\033[38;2;60;86;127mr\033[38;2;58;84;125mj\033[38;2;59;85;125mj\033[38;2;54;80;117mf\033[38;2;55;79;118mf\033[38;2;58;82;122mj\033[38;2;56;82;122mjj\033[38;2;57;82;121mjj\033[38;2;56;80;120mf\033[38;2;56;78;118mf\033[38;2;57;76;117mf\033[38;2;56;78;115mf\033[38;2;54;77;112mf\033[38;2;55;76;111mt\033[38;2;45;65;97m?\033[38;2;47;66;99m?\033[38;2;50;72;107m1\033[38;2;54;79;112mf\033[38;2;52;73;104m1\033[38;2;44;50;66m~\033[38;2;158;151;140mQ\033[38;2;214;198;171mk\033[38;2;231;211;178ma\033[38;2;209;191;163md\033[38;2;195;179;157mq\033[38;2;194;180;161mq\033[38;2;196;182;162mp\033[38;2;198;184;163mp\033[38;2;199;185;162mp\033[38;2;204;189;166md\033[38;2;186;174;155mw\033[38;2;87;91;95mr\033[38;2;159;147;126mL\033[38;2;183;176;157mw\033[38;2;53;67;94m?\033[38;2;48;65;87m-\033[38;2;29;38;55ml\033[38;2;29;37;55mll\033[38;2;24;33;50mI\033[38;2;45;47;53mi\033[38;2;52;52;57m~\033[38;2;24;33;51ml\033[38;2;26;37;54ml\033[38;2;27;36;53ml\033[38;2;24;33;50mI\033[38;2;22;29;48mI\033[38;2;31;45;64mi\033[38;2;40;59;74m+\033[38;2;42;62;79m_\033[38;2;50;68;84m-\033[38;2;178;183;189mp\033[38;2;255;255;255m$$\033[0m                 \033[0m");
  $display("\033[0m      \033[38;2;255;0;0mfff\033[0m        \033[38;2;255;255;255m$\033[38;2;247;248;248mB\033[38;2;134;149;171mQ\033[38;2;77;101;137mu\033[38;2;168;180;196mp\033[38;2;255;255;255m$\033[38;2;157;171;188mw\033[38;2;56;81;120mf\033[38;2;61;84;125mr\033[38;2;58;84;124mjj\033[38;2;56;81;117mf\033[38;2;55;81;117mf\033[38;2;57;83;123mj\033[38;2;56;82;122mjj\033[38;2;56;81;120mf\033[38;2;53;76;114mf\033[38;2;57;80;117mf\033[38;2;56;78;117mf\033[38;2;56;75;116mf\033[38;2;58;75;117mf\033[38;2;58;77;116mf\033[38;2;53;73;107mt\033[38;2;52;75;107mt\033[38;2;53;76;110mt\033[38;2;70;81;105mf\033[38;2;82;92;107mr\033[38;2;49;70;101m1\033[38;2;65;79;102mf\033[38;2;103;98;90mx\033[38;2;252;234;195mW\033[38;2;253;232;192mW\033[38;2;247;227;189mM\033[38;2;246;226;189m#\033[38;2;241;222;187m#\033[38;2;233;214;182mo\033[38;2;225;207;178ma\033[38;2;217;202;173mk\033[38;2;213;197;169mb\033[38;2;217;200;174mk\033[38;2;233;216;186mo\033[38;2;223;212;181ma\033[38;2;136;130;114mY\033[38;2;191;180;157mq\033[38;2;109;111;118mv\033[38;2;39;53;77m+\033[38;2;30;39;57m!\033[38;2;29;37;56ml\033[38;2;28;36;55ml\033[38;2;30;37;51ml\033[38;2;62;57;50m+\033[38;2;118;103;85mn\033[38;2;23;28;44m;\033[38;2;27;35;53ml\033[38;2;27;34;53ml\033[38;2;25;33;51ml\033[38;2;24;29;48mI\033[38;2;27;38;55ml\033[38;2;39;58;72m+\033[38;2;44;63;77m_\033[38;2;39;61;72m+\033[38;2;54;70;89m?\033[38;2;126;136;152mJ\033[38;2;167;174;184mw\033[38;2;199;204;209ma\033[38;2;216;218;223m#\033[38;2;214;217;222m#\033[38;2;202;206;212ma\033[38;2;241;242;244m%%\033[38;2;255;255;255m$\033[0m           \033[0m");
  $display("\033[0m                \033[38;2;255;255;255m$\033[38;2;238;239;240m%%\033[38;2;109;128;155mY\033[38;2;106;127;157mY\033[38;2;214;220;229mM\033[38;2;255;255;255m$\033[38;2;181;190;206mb\033[38;2;61;85;124mr\033[38;2;58;83;123mj\033[38;2;58;84;124mj\033[38;2;57;84;124mj\033[38;2;55;82;120mf\033[38;2;55;80;115mf\033[38;2;58;83;122mj\033[38;2;57;82;122mj\033[38;2;56;82;122mj\033[38;2;56;82;121mj\033[38;2;52;76;112mt\033[38;2;53;75;108mt\033[38;2;56;78;116mf\033[38;2;57;76;118mf\033[38;2;58;75;118mf\033[38;2;57;77;115mf\033[38;2;56;78;113mf\033[38;2;50;72;106m1\033[38;2;54;77;109mt\033[38;2;49;71;102m1\033[38;2;156;151;143mQ\033[38;2;243;226;192m#\033[38;2;190;176;158mw\033[38;2;181;171;153mm\033[38;2;199;183;157mq\033[38;2;223;206;174mh\033[38;2;227;209;176ma\033[38;2;231;212;179mo\033[38;2;235;215;183mo\033[38;2;237;217;185m*\033[38;2;236;217;184m*\033[38;2;232;215;183mo\033[38;2;234;218;184m*\033[38;2;244;226;193mM\033[38;2;246;226;193mM\033[38;2;246;224;189m#\033[38;2;247;226;190mM\033[38;2;243;225;190m#\033[38;2;222;206;177mh\033[38;2;169;159;144m0\033[38;2;42;47;61m~\033[38;2;27;34;49ml\033[38;2;37;43;55mi\033[38;2;27;30;43mI\033[38;2;92;82;78mf\033[38;2;93;80;63mt\033[38;2;158;137;105mU\033[38;2;43;42;48m!\033[38;2;26;33;50ml\033[38;2;26;37;54ml\033[38;2;25;33;51ml\033[38;2;25;29;47mI\033[38;2;25;35;52ml\033[38;2;34;54;68m~\033[38;2;38;60;76m+\033[38;2;38;60;78m+\033[38;2;79;90;100mj\033[38;2;210;213;215m*\033[38;2;145;154;166m0\033[38;2;127;138;153mJ\033[38;2;141;151;165mQ\033[38;2;152;160;172mO\033[38;2;175;181;190mp\033[38;2;237;239;240m8\033[38;2;255;255;255m$\033[0m           \033[0m");
  $display("\033[0m               \033[38;2;255;255;255m$\033[38;2;237;238;238m8\033[38;2;99;119;147mz\033[38;2;122;141;168mC\033[38;2;243;244;246mB\033[38;2;255;255;255m$\033[38;2;214;217;226m#\033[38;2;76;100;138mu\033[38;2;57;80;123mj\033[38;2;57;84;124mj\033[38;2;56;86;124mj\033[38;2;56;82;121mj\033[38;2;53;78;116mf\033[38;2;57;83;122mj\033[38;2;56;82;122mj\033[38;2;57;82;122mjj\033[38;2;57;81;118mf\033[38;2;50;73;106m1\033[38;2;57;78;114mf\033[38;2;56;76;117mf\033[38;2;56;75;117mff\033[38;2;53;75;113mt\033[38;2;54;77;109mt\033[38;2;52;74;109mt\033[38;2;52;75;110mt\033[38;2;51;70;97m1\033[38;2;198;186;165mp\033[38;2;252;232;195mW\033[38;2;253;231;194mW\033[38;2;245;225;189m#\033[38;2;157;140;119mJ\033[38;2;126;112;100mv\033[38;2;126;118;107mz\033[38;2;132;127;117mX\033[38;2;165;158;147m0\033[38;2;129;121;111mz\033[38;2;118;109;97mv\033[38;2;112;100;86mn\033[38;2;150;134;118mU\033[38;2;240;223;195m#\033[38;2;242;225;195m#\033[38;2;242;224;191m###\033[38;2;246;227;194mM\033[38;2;237;218;184m*\033[38;2;187;166;134mZ\033[38;2;148;129;102mY\033[38;2;160;139;109mJ\033[38;2;148;124;96mX\033[38;2;122;103;84mn\033[38;2;116;98;78mx\033[38;2;166;143;107mJ\033[38;2;66;62;57m_\033[38;2;22;30;47mI\033[38;2;28;36;52ml\033[38;2;25;30;47mI\033[38;2;27;31;48mI\033[38;2;25;34;50ml\033[38;2;31;46;60mi\033[38;2;37;56;71m+\033[38;2;42;63;80m_\033[38;2;35;52;70m~\033[38;2;172;174;175mw\033[38;2;255;255;255m$$$$$\033[0m             \033[0m");
  $display("\033[0m              \033[38;2;255;255;255m$\033[38;2;241;241;241m%%\033[38;2;102;120;146mX\033[38;2;118;137;165mC\033[38;2;249;251;251m@\033[0m \033[38;2;255;255;255m$\033[38;2;138;153;177m0\033[38;2;49;75;116mt\033[38;2;60;84;125mj\033[38;2;57;84;124mj\033[38;2;56;85;122mj\033[38;2;52;77;114mf\033[38;2;57;84;122mj\033[38;2;56;84;123mj\033[38;2;56;82;122mj\033[38;2;57;82;122mjj\033[38;2;53;77;113mf\033[38;2;51;74;107mt\033[38;2;56;78;116mf\033[38;2;54;76;116mf\033[38;2;54;76;112mt\033[38;2;55;76;116mf\033[38;2;49;68;101m1\033[38;2;50;72;101m1\033[38;2;53;77;111mt\033[38;2;49;73;107m1\033[38;2;54;70;101m1\033[38;2;205;191;171mb\033[38;2;250;229;194mM\033[38;2;244;225;190m#\033[38;2;244;225;188m#\033[38;2;247;227;189mM\033[38;2;243;231;197mM\033[38;2;236;235;220m&\033[38;2;231;234;220mW\033[38;2;230;232;217mW\033[38;2;229;230;220mW\033[38;2;228;225;206m#\033[38;2;232;215;184mo\033[38;2;231;215;182mo\033[38;2;240;224;194m#\033[38;2;242;225;197mM\033[38;2;241;224;195m#\033[38;2;241;224;194m#\033[38;2;239;224;194m#\033[38;2;242;223;191m#\033[38;2;243;225;191m#\033[38;2;239;221;185m*\033[38;2;230;212;177ma\033[38;2;234;217;182mo\033[38;2;187;164;124mO\033[38;2;167;142;107mJ\033[38;2;170;145;112mC\033[38;2;175;148;110mL\033[38;2;74;65;60m-\033[38;2;24;28;46mI\033[38;2;30;32;49ml\033[38;2;24;30;46mI\033[38;2;24;34;50ml\033[38;2;23;33;50mI\033[38;2;26;40;56ml\033[38;2;31;50;64mi\033[38;2;44;63;79m_\033[38;2;39;58;78m+\033[38;2;89;96;107mx\033[38;2;247;245;243mB\033[0m                 \033[0m");
  $display("\033[0m             \033[38;2;255;255;255m$\033[38;2;255;255;252m$\033[38;2;125;141;164mC\033[38;2;86;109;143mv\033[38;2;234;237;241m8\033[38;2;255;255;255m$\033[0m \033[38;2;244;244;247mB\033[38;2;94;115;146mz\033[38;2;55;81;120mf\033[38;2;59;84;124mj\033[38;2;59;85;124mj\033[38;2;54;80;114mf\033[38;2;55;80;118mf\033[38;2;57;85;125mj\033[38;2;55;83;122mj\033[38;2;56;82;122mj\033[38;2;57;82;122mj\033[38;2;56;81;121mj\033[38;2;49;73;109mt\033[38;2;54;77;112mf\033[38;2;54;77;114mf\033[38;2;54;76;113mf\033[38;2;54;76;111mt\033[38;2;55;77;114mf\033[38;2;44;61;88m-\033[38;2;45;63;91m-\033[38;2;55;80;112mf\033[38;2;49;73;106m1\033[38;2;39;60;97m-\033[38;2;161;156;149m0\033[38;2;253;233;198mW\033[38;2;244;226;191m##\033[38;2;244;225;189m#\033[38;2;238;228;199mM\033[38;2;232;232;220mW\033[38;2;230;230;218mW\033[38;2;231;231;219mW\033[38;2;231;233;220mW\033[38;2;238;230;207mW\033[38;2;242;225;190m#\033[38;2;241;225;192m#\033[38;2;241;224;194m####\033[38;2;241;224;195m#\033[38;2;240;223;191m#\033[38;2;244;225;191m#\033[38;2;232;215;185mo\033[38;2;120;106;93mu\033[38;2;130;121;105mz\033[38;2;156;141;116mJ\033[38;2;152;128;98mY\033[38;2;171;146;111mC\033[38;2;177;147;110mL\033[38;2;99;85;74mj\033[38;2;28;30;46mI\033[38;2;26;30;48mI\033[38;2;28;33;49ml\033[38;2;26;34;51ml\033[38;2;25;33;50ml\033[38;2;25;35;51ml\033[38;2;29;45;61mi\033[38;2;43;62;80m_\033[38;2;41;62;81m_\033[38;2;40;57;75m+\033[38;2;198;198;198mh\033[38;2;255;255;255m$\033[0m                \033[0m");
  $display("\033[0m             \033[38;2;255;255;255m$\033[38;2;182;189;199mb\033[38;2;58;83;121mj\033[38;2;200;208;219mo\033[38;2;255;255;255m$\033[0m \033[38;2;255;255;255m$\033[38;2;220;222;230mM\033[38;2;68;90;128mx\033[38;2;58;84;122mj\033[38;2;60;86;123mj\033[38;2;58;83;120mj\033[38;2;54;77;114mf\033[38;2;58;84;123mj\033[38;2;56;84;123mj\033[38;2;55;83;122mj\033[38;2;56;82;120mjj\033[38;2;55;81;118mf\033[38;2;48;72;106m1\033[38;2;55;76;114mf\033[38;2;55;75;114mf\033[38;2;55;77;114mf\033[38;2;54;77;113mf\033[38;2;55;78;113mf\033[38;2;42;59;85m_\033[38;2;37;50;72m~\033[38;2;55;79;111mf\033[38;2;56;76;104mt\033[38;2;125;131;137mU\033[38;2;83;91;104mr\033[38;2;223;209;184ma\033[38;2;249;232;198mW\033[38;2;242;226;192m#\033[38;2;242;225;189m#\033[38;2;236;230;204mM\033[38;2;232;232;220mW\033[38;2;232;232;219mW\033[38;2;231;233;220mW\033[38;2;232;233;218mW\033[38;2;239;226;198mM\033[38;2;241;224;194m##\033[38;2;240;223;193m#\033[38;2;240;223;192m#\033[38;2;240;223;191m#\033[38;2;241;224;192m#\033[38;2;240;224;192m#\033[38;2;241;225;194m#\033[38;2;240;226;194m#\033[38;2;242;225;189m#\033[38;2;237;217;182m*\033[38;2;202;189;162mp\033[38;2;137;136;120mU\033[38;2;76;72;64m?\033[38;2;113;98;79mx\033[38;2;168;145;106mJ\033[38;2;92;84;72mf\033[38;2;28;31;45mI\033[38;2;30;33;51ml\033[38;2;32;35;52ml\033[38;2;29;31;49ml\033[38;2;24;29;46mI\033[38;2;25;30;46mI\033[38;2;29;42;57m!\033[38;2;41;59;80m_\033[38;2;36;56;76m+\033[38;2;32;52;73m~\033[38;2;137;140;145mC\033[38;2;255;255;255m$\033[0m                \033[0m");
  $display("\033[0m            \033[38;2;255;255;255m$\033[38;2;248;248;247mB\033[38;2;90;110;138mv\033[38;2;92;115;148mz\033[38;2;250;250;251m@\033[0m  \033[38;2;255;255;255m$\033[38;2;179;186;200md\033[38;2;53;78;118mf\033[38;2;59;86;123mj\033[38;2;59;86;122mj\033[38;2;54;77;116mf\033[38;2;58;80;120mj\033[38;2;57;84;124mj\033[38;2;54;83;122mj\033[38;2;55;83;122mj\033[38;2;55;82;120mff\033[38;2;53;78;114mf\033[38;2;49;71;105m1\033[38;2;56;75;117mf\033[38;2;56;74;115mf\033[38;2;55;75;114mf\033[38;2;53;76;110mt\033[38;2;53;78;111mt\033[38;2;43;61;89m-\033[38;2;30;40;58m!\033[38;2;50;67;102m1\033[38;2;65;78;102mf\033[38;2;231;216;188mo\033[38;2;194;182;162mq\033[38;2;133;128;122mY\033[38;2;209;195;169mb\033[38;2;238;223;190m#\033[38;2;240;224;188m#\033[38;2;235;232;209mW\033[38;2;231;233;220mW\033[38;2;231;232;220mW\033[38;2;231;234;218mW\033[38;2;234;231;215mW\033[38;2;241;225;193m#\033[38;2;242;224;192m#\033[38;2;242;224;195m#\033[38;2;241;224;195m#\033[38;2;240;224;193m#\033[38;2;240;224;192m#\033[38;2;240;224;191m##\033[38;2;241;224;194m#\033[38;2;239;221;188m#\033[38;2;241;222;189m#\033[38;2;244;225;187m#\033[38;2;244;229;198mM\033[38;2;198;196;175mb\033[38;2;169;167;146mO\033[38;2;164;149;119mL\033[38;2;105;91;76mr\033[38;2;22;30;46mI\033[38;2;29;35;52ml\033[38;2;32;34;52ml\033[38;2;30;33;50ml\033[38;2;26;29;46mI\033[38;2;25;28;45mI\033[38;2;28;31;48mI\033[38;2;29;40;55m!\033[38;2;39;58;79m+\033[38;2;36;56;73m+\033[38;2;30;50;71m~\033[38;2;114;121;131mX\033[38;2;255;255;255m$\033[0m                \033[0m");
  $display("\033[0m            \033[38;2;255;255;255m$\033[38;2;238;238;239m8\033[38;2;76;98;130mn\033[38;2;75;100;135mn\033[38;2;231;233;238m8\033[38;2;255;255;255m$\033[0m \033[38;2;255;255;255m$\033[38;2;141;152;174m0\033[38;2;51;76;115mt\033[38;2;58;85;122mj\033[38;2;57;81;119mf\033[38;2;52;77;116mf\033[38;2;56;83;123mj\033[38;2;55;83;122mjj\033[38;2;55;82;122mj\033[38;2;54;81;121mf\033[38;2;52;81;120mf\033[38;2;47;70;102m1\033[38;2;51;69;103m1\033[38;2;57;74;117mf\033[38;2;56;73;116mf\033[38;2;56;73;115mf\033[38;2;54;74;111mt\033[38;2;52;76;111mt\033[38;2;50;68;101m1\033[38;2;29;39;60m!\033[38;2;37;52;78m+\033[38;2;66;77;96mt\033[38;2;220;203;176mh\033[38;2;255;235;198mW\033[38;2;235;215;185mo\033[38;2;202;186;162mp\033[38;2;216;202;172mk\033[38;2;230;214;182mo\033[38;2;233;231;213mW\033[38;2;231;234;221mW\033[38;2;230;232;221mW\033[38;2;230;233;220mW\033[38;2;236;229;210mW\033[38;2;240;224;189m#\033[38;2;241;224;192m#\033[38;2;241;224;195m#\033[38;2;240;223;195m#\033[38;2;240;223;193m##\033[38;2;240;223;191m#\033[38;2;239;223;190m#\033[38;2;240;223;190m#\033[38;2;242;223;190m##\033[38;2;239;222;188m#\033[38;2;237;228;207mM\033[38;2;204;203;188mh\033[38;2;171;162;137m0\033[38;2;163;143;111mJ\033[38;2;48;46;52mi\033[38;2;28;33;51ml\033[38;2;32;35;54ml\033[38;2;29;33;51ml\033[38;2;23;30;46mI\033[38;2;23;29;46mI\033[38;2;24;32;49mI\033[38;2;25;32;49mI\033[38;2;26;39;53ml\033[38;2;40;60;76m+\033[38;2;39;58;75m+\033[38;2;34;54;68m~\033[38;2;173;176;178mw\033[38;2;255;255;255m$\033[0m                \033[0m");
  $display("\033[0m             \033[38;2;255;255;255m$\033[38;2;148;161;178mZ\033[38;2;42;70;111m1\033[38;2;133;150;173mQ\033[38;2;255;255;255m$$$\033[38;2;165;175;192mq\033[38;2;50;76;113mt\033[38;2;59;83;120mj\033[38;2;54;77;114mf\033[38;2;55;81;120mf\033[38;2;54;83;122mj\033[38;2;55;82;121mj\033[38;2;55;83;121mj\033[38;2;55;81;120mf\033[38;2;54;80;120mf\033[38;2;52;81;118mf\033[38;2;40;57;82m_\033[38;2;50;71;105m1\033[38;2;56;74;116mf\033[38;2;56;73;116mf\033[38;2;56;73;115mf\033[38;2;54;74;110mt\033[38;2;53;76;109mt\033[38;2;54;74;108mt\033[38;2;36;47;70m~\033[38;2;29;41;61m!\033[38;2;59;67;81m?\033[38;2;198;175;145mw\033[38;2;248;232;195mW\033[38;2;244;228;191mM\033[38;2;247;229;192mM\033[38;2;244;225;188m#\033[38;2;240;227;197mM\033[38;2;232;233;220mW\033[38;2;231;233;220mWW\033[38;2;231;234;219mW\033[38;2;238;228;204mM\033[38;2;241;224;189m#\033[38;2;241;225;193m#\033[38;2;243;226;196mM\033[38;2;243;227;196mM\033[38;2;241;226;192m#\033[38;2;239;223;191m#\033[38;2;242;227;194mM\033[38;2;242;226;192m#\033[38;2;239;222;189m#\033[38;2;240;222;189m#\033[38;2;240;221;187m#\033[38;2;236;222;190m#\033[38;2;235;230;216mW\033[38;2;191;189;170mp\033[38;2;173;160;126m0\033[38;2;125;110;92mv\033[38;2;27;31;48mI\033[38;2;32;34;53ml\033[38;2;30;34;53ml\033[38;2;27;34;52ml\033[38;2;24;33;49mI\033[38;2;25;34;50ml\033[38;2;26;35;52ml\033[38;2;25;33;50ml\033[38;2;27;40;55ml\033[38;2;39;60;75m+\033[38;2;34;54;75m+\033[38;2;82;94;106mr\033[38;2;250;248;247m@\033[38;2;255;255;255m$\033[0m                \033[0m");
  $display("\033[0m             \033[38;2;255;255;255m$\033[38;2;240;240;241m%%\033[38;2;130;146;168mL\033[38;2;51;78;116mf\033[38;2;108;127;156mY\033[38;2;175;186;201md\033[38;2;207;214;223m*\033[38;2;178;187;201md\033[38;2;58;79;115mf\033[38;2;60;80;116mf\033[38;2;52;75;111mt\033[38;2;56;82;122mj\033[38;2;55;83;122mj\033[38;2;55;82;120mf\033[38;2;56;82;119mff\033[38;2;55;82;119mf\033[38;2;51;76;109mt\033[38;2;34;47;68mi\033[38;2;52;72;107mt\033[38;2;55;74;117mf\033[38;2;55;74;116mf\033[38;2;55;74;115mf\033[38;2;54;74;112mt\033[38;2;53;75;109mt\033[38;2;53;76;111mt\033[38;2;43;61;89m-\033[38;2;27;39;57m!\033[38;2;38;48;64m~\033[38;2;140;120;100mz\033[38;2;218;195;160mb\033[38;2;245;230;196mM\033[38;2;244;227;189m#\033[38;2;242;225;188m#\033[38;2;236;229;205mM\033[38;2;232;233;222mW\033[38;2;231;232;219mW\033[38;2;230;232;219mW\033[38;2;231;233;217mW\033[38;2;240;225;194m#\033[38;2;244;224;189m#\033[38;2;240;222;191m#\033[38;2;220;197;171mk\033[38;2;197;165;141mm\033[38;2;177;140;116mL\033[38;2;160;124;106mY\033[38;2;134;110;95mc\033[38;2;213;196;170mb\033[38;2;245;226;192mM\033[38;2;239;223;189m#\033[38;2;238;223;186m*\033[38;2;237;228;203mM\033[38;2;207;207;189mh\033[38;2;174;166;139mO\033[38;2;165;148;113mC\033[38;2;59;54;54m+\033[38;2;24;30;50mI\033[38;2;29;36;54ml\033[38;2;26;35;52ml\033[38;2;25;33;51ml\033[38;2;26;31;50mI\033[38;2;26;33;51ml\033[38;2;26;35;52ml\033[38;2;25;33;50ml\033[38;2;29;42;58m!\033[38;2;40;61;77m_\033[38;2;35;57;75m+\033[38;2;33;53;69m~\033[38;2;182;187;192md\033[38;2;255;255;255m$\033[0m                \033[0m");
  $display("\033[0m              \033[38;2;255;255;255m$\033[38;2;255;255;253m$\033[38;2;179;186;196md\033[38;2;103;122;148mX\033[38;2;72;96;130mn\033[38;2;73;98;132mn\033[38;2;66;91;125mr\033[38;2;59;82;115mf\033[38;2;56;79;112mf\033[38;2;52;74;110mt\033[38;2;57;82;122mj\033[38;2;56;81;121mj\033[38;2;56;82;119mff\033[38;2;55;81;118mf\033[38;2;56;81;120mf\033[38;2;44;66;94m?\033[38;2;33;43;65mi\033[38;2;54;72;109mt\033[38;2;55;74;117mf\033[38;2;55;74;116mf\033[38;2;55;74;115mf\033[38;2;54;74;112mt\033[38;2;51;73;108mt\033[38;2;52;75;110mt\033[38;2;51;72;103m1\033[38;2;34;44;62mi\033[38;2;31;40;53m!\033[38;2;28;36;47ml\033[38;2;125;107;88mu\033[38;2;200;178;145mw\033[38;2;232;213;179mo\033[38;2;244;226;190m#\033[38;2;239;232;207mW\033[38;2;234;234;222m&\033[38;2;231;232;220mW\033[38;2;230;232;220mW\033[38;2;231;233;214mW\033[38;2;241;225;191m#\033[38;2;244;223;189m#\033[38;2;192;156;132mO\033[38;2;177;127;110mJ\033[38;2;183;127;113mC\033[38;2;183;126;111mC\033[38;2;177;121;105mU\033[38;2;132;85;73mx\033[38;2;165;146;125mL\033[38;2;248;229;192mM\033[38;2;243;225;189m#\033[38;2;235;220;186m*\033[38;2;202;195;174mb\033[38;2;179;174;151mm\033[38;2;169;156;129mQ\033[38;2;86;77;73mt\033[38;2;24;29;46mI\033[38;2;30;35;52ml\033[38;2;29;35;53ml\033[38;2;27;35;53ml\033[38;2;25;31;48mI\033[38;2;26;31;50mI\033[38;2;26;33;51ml\033[38;2;26;35;52ml\033[38;2;25;32;50mI\033[38;2;31;46;62mi\033[38;2;37;56;75m+\033[38;2;64;80;95mt\033[38;2;108;123;134mz\033[38;2;72;89;103mj\033[38;2;240;240;240m%%\033[38;2;255;255;255m$\033[0m               \033[0m");
  $display("\033[0m                \033[38;2;255;255;255m$\033[38;2;252;250;247m@\033[38;2;200;204;207ma\033[38;2;171;178;184mq\033[38;2;177;185;189mp\033[38;2;199;202;208ma\033[38;2;74;93;123mx\033[38;2;50;72;110mt\033[38;2;57;83;121mj\033[38;2;57;83;120mj\033[38;2;56;83;118mf\033[38;2;55;82;118mf\033[38;2;54;80;117mf\033[38;2;55;81;118mf\033[38;2;41;58;85m_\033[38;2;32;44;63mi\033[38;2;53;72;108mt\033[38;2;53;74;114mt\033[38;2;54;74;115mf\033[38;2;54;73;115mt\033[38;2;54;74;111mt\033[38;2;51;74;108mtt\033[38;2;53;74;107mt\033[38;2;37;50;73m~\033[38;2;32;39;54m!\033[38;2;21;30;48mI\033[38;2;116;102;84mn\033[38;2;182;156;119mQ\033[38;2;181;153;119mQ\033[38;2;195;171;134mZ\033[38;2;211;196;167mb\033[38;2;225;221;205m#\033[38;2;232;234;223mW\033[38;2;232;237;225m&\033[38;2;236;233;212mW\033[38;2;244;224;188m#\033[38;2;244;224;189m#\033[38;2;235;213;180mo\033[38;2;235;209;177mo\033[38;2;237;208;177mo\033[38;2;233;201;172mh\033[38;2;225;191;163mb\033[38;2;219;189;160mb\033[38;2;233;211;178mo\033[38;2;242;221;183m*\033[38;2;217;200;168mk\033[38;2;190;179;156mw\033[38;2;170;166;147mO\033[38;2;135;133;120mY\033[38;2;63;63;64m-\033[38;2;26;29;49mI\033[38;2;31;34;54ml\033[38;2;29;32;51ml\033[38;2;28;34;52ml\033[38;2;26;32;50ml\033[38;2;25;30;47mI\033[38;2;26;33;51ml\033[38;2;25;34;52ml\033[38;2;26;35;52ml\033[38;2;25;33;48mI\033[38;2;34;52;68m~\033[38;2;29;50;70mi\033[38;2;155;161;167mO\033[38;2;255;255;255m$\033[38;2;78;91;110mr\033[38;2;164;169;178mm\033[38;2;255;255;255m$\033[0m               \033[0m");
  $display("\033[0m                     \033[38;2;255;255;255m$\033[38;2;177;185;191mp\033[38;2;54;75;107mt\033[38;2;58;82;117mf\033[38;2;58;82;119mj\033[38;2;58;81;117mff\033[38;2;57;80;117mf\033[38;2;57;79;114mf\033[38;2;39;53;78m+\033[38;2;32;44;61mi\033[38;2;50;69;104m1\033[38;2;53;76;110mt\033[38;2;53;75;112mt\033[38;2;55;73;114mt\033[38;2;55;75;111mt\033[38;2;53;76;110mt\033[38;2;52;75;109mt\033[38;2;53;76;110mt\033[38;2;43;59;84m_\033[38;2;30;36;52ml\033[38;2;37;37;51m!\033[38;2;150;129;103mY\033[38;2;184;156;118mQ\033[38;2;181;154;117mQ\033[38;2;179;153;115mQ\033[38;2;178;151;115mL\033[38;2;182;156;121m0\033[38;2;192;173;144mm\033[38;2;204;197;175mb\033[38;2;224;217;193mo\033[38;2;242;225;191m#\033[38;2;251;232;193mW\033[38;2;251;230;193mM\033[38;2;246;226;190m#\033[38;2;244;225;189m#\033[38;2;247;228;191mM\033[38;2;252;232;194mW\033[38;2;249;225;189mM\033[38;2;223;197;163mk\033[38;2;183;162;132mO\033[38;2;148;142;122mJ\033[38;2;111;109;104mv\033[38;2;62;64;71m-\033[38;2;28;34;50ml\033[38;2;25;33;52ml\033[38;2;28;34;53ml\033[38;2;29;34;53ml\033[38;2;26;31;50mI\033[38;2;27;34;52ml\033[38;2;24;31;49mI\033[38;2;25;33;50ml\033[38;2;26;35;52mll\033[38;2;26;34;52ml\033[38;2;27;38;53ml\033[38;2;28;47;66mi\033[38;2;125;136;148mJ\033[38;2;255;255;255m$$\033[38;2;165;171;183mw\033[38;2;94;103;123mu\033[38;2;255;255;255m$$\033[0m              \033[0m");
  $display("\033[0m                     \033[38;2;255;255;255m$\033[38;2;227;229;230mW\033[38;2;64;86;116mj\033[38;2;50;71;102m1\033[38;2;58;80;114mf\033[38;2;57;81;114mf\033[38;2;57;79;113mf\033[38;2;56;80;115mf\033[38;2;57;79;112mf\033[38;2;40;53;76m+\033[38;2;36;42;63mi\033[38;2;48;66;100m?\033[38;2;53;76;113mt\033[38;2;54;74;113mt\033[38;2;54;74;111mt\033[38;2;54;75;110mt\033[38;2;53;75;110mt\033[38;2;53;75;109mt\033[38;2;53;76;109mt\033[38;2;48;68;98m?\033[38;2;31;37;57m!\033[38;2;42;43;57mi\033[38;2;151;147;134mL\033[38;2;164;147;121mL\033[38;2;173;148;112mL\033[38;2;180;152;115mQ\033[38;2;181;154;116mQ\033[38;2;182;153;115mQ\033[38;2;181;152;112mL\033[38;2;178;150;111mL\033[38;2;180;155;118mQ\033[38;2;158;143;118mJ\033[38;2;136;129;117mY\033[38;2;192;176;155mw\033[38;2;228;210;180ma\033[38;2;242;222;188m#\033[38;2;221;203;171mh\033[38;2;183;165;140mZ\033[38;2;133;117;102mz\033[38;2;86;78;75mt\033[38;2;55;57;63m+\033[38;2;34;42;56m!\033[38;2;23;33;48mI\033[38;2;24;34;52ml\033[38;2;28;37;55ml\033[38;2;28;37;54ml\033[38;2;26;34;52ml\033[38;2;27;34;52ml\033[38;2;24;31;49mI\033[38;2;26;33;51ml\033[38;2;24;31;49mI\033[38;2;25;34;51ml\033[38;2;25;35;52ml\033[38;2;26;34;52ml\033[38;2;24;33;51ml\033[38;2;23;40;57ml\033[38;2;108;122;134mz\033[38;2;240;242;242m%%\033[38;2;255;255;255m$$\033[38;2;216;218;223m#\033[38;2;84;95;118mn\033[38;2;245;245;247mB\033[38;2;255;255;255m$\033[0m              \033[0m");
  $display("\033[0m                \033[38;2;251;251;251m@\033[38;2;255;255;255m$$\033[0m \033[38;2;255;255;255m$$\033[38;2;150;163;182mZ\033[38;2;62;87;122mr\033[38;2;53;75;103mt\033[38;2;41;58;85m_\033[38;2;48;68;103m1\033[38;2;57;80;116mf\033[38;2;57;80;113mf\033[38;2;57;79;114mf\033[38;2;42;55;80m_\033[38;2;37;42;61mi\033[38;2;44;59;85m_\033[38;2;54;77;114mf\033[38;2;53;75;113mt\033[38;2;53;75;112mt\033[38;2;53;76;110mt\033[38;2;52;74;109mt\033[38;2;52;75;109mt\033[38;2;51;74;108mt\033[38;2;51;73;107mt\033[38;2;39;51;77m+\033[38;2;25;31;49mI\033[38;2;122;128;129mY\033[38;2;170;176;163mm\033[38;2;159;157;142mQ\033[38;2;161;146;123mC\033[38;2;171;147;113mC\033[38;2;180;151;112mL\033[38;2;181;154;114mQ\033[38;2;182;153;114mQ\033[38;2;180;152;113mL\033[38;2;103;95;88mx\033[38;2;21;28;47mI\033[38;2;34;40;57m!\033[38;2;56;62;71m-\033[38;2;71;75;82m1\033[38;2;48;53;61m+\033[38;2;30;39;52ml\033[38;2;24;35;51ml\033[38;2;25;35;53ml\033[38;2;29;37;56ml\033[38;2;30;37;55ml\033[38;2;29;38;52ml\033[38;2;29;37;55ml\033[38;2;29;38;55ml\033[38;2;26;35;52ml\033[38;2;26;34;51ml\033[38;2;27;34;52ml\033[38;2;23;30;48mI\033[38;2;26;33;51ml\033[38;2;26;35;52mll\033[38;2;26;34;52ml\033[38;2;24;32;48mI\033[38;2;20;31;49mI\033[38;2;95;108;123mv\033[38;2;241;242;242m%%\033[38;2;255;255;255m$\033[0m \033[38;2;255;255;255m$\033[38;2;173;179;189mp\033[38;2;109;118;137mz\033[38;2;255;255;255m$$\033[0m              \033[0m");
  $display("\033[0m               \033[38;2;255;255;255m$$\033[38;2;241;244;248mB\033[38;2;202;209;219mo\033[38;2;191;200;211mh\033[38;2;184;192;206mk\033[38;2;152;167;189mm\033[38;2;142;157;178mO\033[38;2;174;184;199md\033[38;2;56;81;116mf\033[38;2;110;122;133mz\033[38;2;105;113;121mc\033[38;2;46;62;88m-\033[38;2;54;76;107mt\033[38;2;57;82;115mf\033[38;2;47;60;87m-\033[38;2;39;45;62mi\033[38;2;39;53;72m+\033[38;2;54;76;112mt\033[38;2;53;76;112mt\033[38;2;53;77;111mt\033[38;2;53;76;110mt\033[38;2;53;76;109mtt\033[38;2;51;74;108mt\033[38;2;51;74;109mt\033[38;2;47;67;98m?\033[38;2;27;36;57ml\033[38;2;54;59;70m_\033[38;2;161;165;155mO\033[38;2;171;175;165mm\033[38;2;166;169;161mZ\033[38;2;160;159;147m0\033[38;2;160;147;125mL\033[38;2;169;146;112mC\033[38;2;179;150;109mL\033[38;2;164;141;109mJ\033[38;2;157;160;150m0\033[38;2;98;102;102mn\033[38;2;27;36;52ml\033[38;2;31;40;59m!\033[38;2;30;40;58m!\033[38;2;31;41;59m!\033[38;2;31;39;57m!\033[38;2;30;37;55ml\033[38;2;29;36;54ml\033[38;2;32;38;57m!\033[38;2;30;37;54ml\033[38;2;29;38;52ml\033[38;2;29;37;56ml\033[38;2;28;37;55ml\033[38;2;25;33;52ml\033[38;2;25;32;51ml\033[38;2;23;30;49mI\033[38;2;23;31;49mI\033[38;2;26;34;52ml\033[38;2;26;35;52mll\033[38;2;25;33;50ml\033[38;2;22;34;50mI\033[38;2;47;62;81m-\033[38;2;213;214;219m*\033[38;2;255;255;255m$\033[0m \033[38;2;255;255;255m$\033[38;2;223;224;228mW\033[38;2;82;93;115mx\033[38;2;212;216;222m#\033[38;2;255;255;255m$\033[0m               \033[0m");
  $display("\033[0m                \033[38;2;255;255;255m$\033[38;2;246;246;250mB\033[38;2;218;222;231mM\033[38;2;200;207;217mo\033[38;2;194;203;214ma\033[38;2;210;216;222m#\033[38;2;255;255;255m$\033[38;2;116;135;163mJ\033[38;2;144;158;175mO\033[38;2;255;255;253m$\033[38;2;255;255;255m$\033[38;2;125;133;140mU\033[38;2;31;44;67mi\033[38;2;45;63;93m-\033[38;2;53;68;98m1\033[38;2;40;46;66m~\033[38;2;37;47;62mi\033[38;2;52;69;100m1\033[38;2;54;77;115mf\033[38;2;53;76;111mt\033[38;2;53;76;110mt\033[38;2;54;77;111mt\033[38;2;53;76;110mt\033[38;2;50;73;107m1\033[38;2;51;72;107m1\033[38;2;52;75;108mt\033[38;2;40;56;84m_\033[38;2;24;32;56ml\033[38;2;76;80;88mf\033[38;2;164;169;156mZ\033[38;2;172;176;160mm\033[38;2;168;172;159mZ\033[38;2;168;171;160mZ\033[38;2;159;159;149m0\033[38;2;156;148;130mL\033[38;2;150;145;128mC\033[38;2;149;153;143mL\033[38;2;167;170;159mZ\033[38;2;81;88;90mj\033[38;2;31;38;55m!\033[38;2;29;37;55ml\033[38;2;33;41;59m!\033[38;2;32;39;58m!\033[38;2;29;36;55ml\033[38;2;29;37;55mll\033[38;2;29;38;54mll\033[38;2;28;38;55ml\033[38;2;28;37;56ml\033[38;2;24;32;51mI\033[38;2;22;29;48mI\033[38;2;24;32;51mI\033[38;2;25;34;51ml\033[38;2;26;35;52ml\033[38;2;25;34;51ml\033[38;2;24;34;51ml\033[38;2;28;40;58m!\033[38;2;27;45;66mi\033[38;2;115;122;130mX\033[38;2;255;255;255m$\033[0m \033[38;2;255;255;255m$\033[38;2;199;203;211ma\033[38;2;94;105;126mv\033[38;2;165;170;182mw\033[38;2;255;255;255m$$\033[0m               \033[0m");
  $display("\033[0m                      \033[38;2;255;255;255m$\033[38;2;129;147;173mQ\033[38;2;181;191;206mb\033[38;2;255;255;255m$\033[38;2;253;252;250m@\033[38;2;146;154;159m0\033[38;2;90;103;117mn\033[38;2;72;79;92mf\033[38;2;37;48;70m~\033[38;2;43;51;73m+\033[38;2;42;48;66m~\033[38;2;45;55;82m_\033[38;2;55;76;114mf\033[38;2;52;76;112mt\033[38;2;54;77;111mtt\033[38;2;53;77;111mt\033[38;2;52;75;107mt\033[38;2;45;64;93m-\033[38;2;47;63;92m-\033[38;2;52;72;106m1\033[38;2;38;52;77m+\033[38;2;26;33;53ml\033[38;2;64;70;79m?\033[38;2;149;152;143mL\033[38;2;172;174;160mm\033[38;2;168;170;156mZ\033[38;2;155;158;149m0\033[38;2;149;155;149mQ\033[38;2;145;152;144mL\033[38;2;151;157;146mQ\033[38;2;163;166;155mO\033[38;2;121;125;118mz\033[38;2;107;115;115mv\033[38;2;65;72;78m?\033[38;2;36;41;56m!\033[38;2;26;33;51ml\033[38;2;26;33;53ml\033[38;2;30;39;57m!\033[38;2;29;38;55mll\033[38;2;29;37;55ml\033[38;2;27;36;53ml\033[38;2;23;32;50mI\033[38;2;23;30;49mI\033[38;2;26;32;50ml\033[38;2;26;35;52ml\033[38;2;25;35;52ml\033[38;2;26;35;52ml\033[38;2;25;34;52ml\033[38;2;26;35;54ml\033[38;2;27;41;56m!\033[38;2;28;48;63mi\033[38;2;145;147;149mL\033[38;2;252;252;253m$\033[38;2;183;187;196md\033[38;2;148;155;169m0\033[38;2;127;136;154mJ\033[38;2;197;201;207mh\033[38;2;255;255;255m$\033[0m                 \033[0m");
  $display("\033[0m                      \033[38;2;255;255;255m$\033[38;2;238;242;245m%%\033[38;2;208;214;221m*\033[38;2;245;244;238m%%\033[38;2;224;223;212m#\033[38;2;210;210;198ma\033[38;2;244;242;229m8\033[38;2;224;223;211m#\033[38;2;90;93;100mr\033[38;2;38;44;67mi\033[38;2;45;52;75m+\033[38;2;42;49;66m~\033[38;2;49;65;91m?\033[38;2;54;79;113mf\033[38;2;54;77;110mt\033[38;2;50;73;108mt\033[38;2;49;73;107m1\033[38;2;53;76;110mt\033[38;2;50;74;106m1\033[38;2;39;54;78m+\033[38;2;39;50;74m+\033[38;2;48;65;94m?\033[38;2;37;49;71m~\033[38;2;29;37;55ml\033[38;2;59;69;81m?\033[38;2;108;117;121mc\033[38;2;138;141;134mJ\033[38;2;165;169;158mZ\033[38;2;156;160;149m0\033[38;2;157;161;150m0\033[38;2;157;162;153m0\033[38;2;133;144;143mC\033[38;2;77;94;112mr\033[38;2;72;99;123mx\033[38;2;109;126;131mX\033[38;2;145;148;142mL\033[38;2;110;114;112mv\033[38;2;53;59;69m_\033[38;2;27;35;54ml\033[38;2;31;40;57m!\033[38;2;30;38;56m!\033[38;2;28;35;53ml\033[38;2;24;31;49mI\033[38;2;25;32;50mI\033[38;2;26;35;52ml\033[38;2;25;35;52mll\033[38;2;26;35;52mlll\033[38;2;24;33;50mI\033[38;2;22;36;51ml\033[38;2;25;47;61m!\033[38;2;105;106;110mu\033[38;2;251;251;250m@\033[38;2;191;194;203mk\033[38;2;198;202;210ma\033[38;2;255;255;255m$$\033[0m                  \033[0m");
  $display("\033[0m                     \033[38;2;255;255;255m$\033[38;2;253;253;250m$\033[38;2;247;245;236m%%\033[38;2;245;243;231m%%\033[38;2;238;237;225m&\033[38;2;239;239;227m8\033[38;2;241;241;228m8\033[38;2;239;238;226m8\033[38;2;244;243;229m8\033[38;2;224;225;215mM\033[38;2;80;84;93mf\033[38;2;42;49;67m~\033[38;2;43;51;70m+\033[38;2;41;49;67m~\033[38;2;48;67;95m?\033[38;2;49;73;107m1\033[38;2;90;103;124mu\033[38;2;80;93;116mx\033[38;2;44;65;100m?\033[38;2;51;74;106mt\033[38;2;53;72;103m1\033[38;2;38;51;71m~\033[38;2;33;43;63mi\033[38;2;43;56;82m_\033[38;2;36;46;67mi\033[38;2;31;40;58m!\033[38;2;55;76;99m1\033[38;2;75;100;122mn\033[38;2;99;118;129mc\033[38;2;118;130;131mY\033[38;2;129;139;139mJ\033[38;2;92;108;119mu\033[38;2;69;95;119mr\033[38;2;73;100;126mn\033[38;2;72;101;126mn\033[38;2;78;100;117mx\033[38;2;159;164;157mO\033[38;2;173;178;164mw\033[38;2;136;141;133mJ\033[38;2;30;39;50ml\033[38;2;30;39;56m!\033[38;2;29;36;54ml\033[38;2;27;34;52ml\033[38;2;27;37;54ml\033[38;2;26;38;54mlll\033[38;2;26;37;53ml\033[38;2;26;35;52ml\033[38;2;27;36;53mll\033[38;2;21;30;47mI\033[38;2;82;88;97mj\033[38;2;89;103;116mn\033[38;2;32;49;65mi\033[38;2;140;153;162mQ\033[38;2;224;229;231mW\033[38;2;212;217;222m#\033[38;2;187;195;201mk\033[38;2;225;229;232mW\033[38;2;255;255;255m$\033[0m                 \033[0m");
  $display("\033[0m                    \033[38;2;255;255;255m$\033[38;2;251;251;249m@\033[38;2;248;248;236mB\033[38;2;237;237;224m&\033[38;2;239;239;227m8\033[38;2;238;238;227m8\033[38;2;237;237;225m&\033[38;2;236;237;223m&\033[38;2;237;238;224m&\033[38;2;238;239;225m8\033[38;2;247;248;232m%%\033[38;2;179;180;175mq\033[38;2;40;44;62mi\033[38;2;50;54;72m+\033[38;2;42;48;65m~\033[38;2;40;51;69m~\033[38;2;40;60;88m_\033[38;2;72;89;112mr\033[38;2;202;205;201mh\033[38;2;96;106;122mv\033[38;2;43;63;94m-\033[38;2;50;69;104m1\033[38;2;50;72;100m1\033[38;2;33;47;67mi\033[38;2;32;42;61mi\033[38;2;42;50;71m+\033[38;2;34;40;58m!\033[38;2;37;47;66m~\033[38;2;70;93;118mr\033[38;2;69;98;124mx\033[38;2;66;92;120mr\033[38;2;60;85;110mf\033[38;2;67;91;115mr\033[38;2;68;90;112mr\033[38;2;74;99;122mx\033[38;2;71;99;124mx\033[38;2;66;93;120mr\033[38;2;107;116;115mv\033[38;2;164;165;150mO\033[38;2;166;168;158mZ\033[38;2;61;68;72m-\033[38;2;25;33;50ml\033[38;2;30;37;55mll\033[38;2;29;38;55mll\033[38;2;27;37;54ml\033[38;2;26;38;54mllll\033[38;2;26;36;54ml\033[38;2;15;23;43m;\033[38;2;121;125;129mX\033[38;2;248;247;247mB\033[38;2;157;165;173mZ\033[38;2;105;123;137mz\033[38;2;123;139;152mJ\033[38;2;137;151;162mQ\033[38;2;145;157;166m0\033[38;2;217;221;225mM\033[38;2;255;255;255m$\033[0m                 \033[0m");
  $display("\033[0m                   \033[38;2;255;255;255m$\033[38;2;252;250;250m@\033[38;2;241;239;227m8\033[38;2;225;225;209m#\033[38;2;228;226;213mM\033[38;2;227;226;215mM\033[38;2;235;235;223m&\033[38;2;237;237;225m&\033[38;2;237;238;224m&\033[38;2;234;235;220mW\033[38;2;233;233;218mW\033[38;2;242;242;230m8\033[38;2;159;159;157mO\033[38;2;55;57;69m_\033[38;2;183;183;181mp\033[38;2;86;92;99mr\033[38;2;26;35;52ml\033[38;2;70;76;88mt\033[38;2;114;125;141mY\033[38;2;124;131;141mU\033[38;2;229;230;218mW\033[38;2;163;167;165mZ\033[38;2;75;85;108mj\033[38;2;44;63;95m-\033[38;2;43;60;88m-\033[38;2;34;43;62mi\033[38;2;35;43;61mi\033[38;2;36;43;62mi\033[38;2;34;38;55m!\033[38;2;49;62;83m-\033[38;2;70;95;120mx\033[38;2;87;105;121mu\033[38;2;119;130;132mY\033[38;2;135;142;137mJ\033[38;2;134;140;132mJ\033[38;2;134;143;138mJ\033[38;2;106;106;83mx\033[38;2;109;105;72mx\033[38;2;123;108;57mx\033[38;2;141;129;84mz\033[38;2;163;164;151mO\033[38;2;133;135;128mU\033[38;2;42;44;57mi\033[38;2;33;36;56m!\033[38;2;31;38;56m!\033[38;2;28;38;53ml\033[38;2;27;38;53ml\033[38;2;29;37;54ml\033[38;2;29;36;54ml\033[38;2;29;37;53ml\033[38;2;27;35;52ml\033[38;2;22;31;48mI\033[38;2;29;36;47ml\033[38;2;27;31;41mI\033[38;2;83;88;90mj\033[38;2;255;255;255m$$$$$$\033[0m                   \033[0m");
  $display("\033[0m                   \033[38;2;255;255;255m$\033[38;2;248;247;242mB\033[38;2;236;236;220m&\033[38;2;237;238;220m&\033[38;2;237;238;222m&\033[38;2;233;233;216mW\033[38;2;223;221;206m#\033[38;2;234;233;220mW\033[38;2;239;240;226m8\033[38;2;234;234;221mW\033[38;2;225;226;213mM\033[38;2;212;212;201mo\033[38;2;161;161;153mO\033[38;2;209;210;198ma\033[38;2;246;246;229m%%\033[38;2;216;217;206m*\033[38;2;109;113;114mv\033[38;2;55;57;69m_\033[38;2;180;180;173mq\033[38;2;169;171;168mm\033[38;2;120;125;129mX\033[38;2;187;190;183md\033[38;2;219;220;207m*\033[38;2;162;166;166mZ\033[38;2;78;93;111mr\033[38;2;39;53;75m+\033[38;2;35;43;60mi\033[38;2;38;43;59mi\033[38;2;40;42;60mi\033[38;2;38;42;53m!\033[38;2;109;102;58mj\033[38;2;140;123;67mv\033[38;2;153;145;106mU\033[38;2;147;147;126mC\033[38;2;152;154;131mL\033[38;2;136;123;81mc\033[38;2;151;125;52mv\033[38;2;154;128;52mv\033[38;2;153;127;53mv\033[38;2;146;120;50mu\033[38;2;139;128;87mz\033[38;2;168;169;156mZ\033[38;2;98;100;100mn\033[38;2;29;30;46mI\033[38;2;37;39;55m!\033[38;2;35;37;53m!\033[38;2;32;36;52ml\033[38;2;32;35;52ml\033[38;2;31;33;51ml\033[38;2;25;28;46mI\033[38;2;34;37;50ml\033[38;2;63;67;66m-\033[38;2;75;79;55m?\033[38;2;24;30;24m,\033[38;2;107;113;106mv\033[38;2;255;255;255m$\033[0m                        \033[0m");
  $display("\033[0m                   \033[38;2;255;255;255m$\033[38;2;252;252;244m@\033[38;2;236;238;222m&\033[38;2;237;238;220m&\033[38;2;236;237;219m&\033[38;2;239;239;220m&\033[38;2;235;233;217mW\033[38;2;191;190;177md\033[38;2;223;224;208m#\033[38;2;237;239;222m&\033[38;2;236;238;222m&\033[38;2;235;237;222m&\033[38;2;241;243;225m8\033[38;2;237;239;222m&\033[38;2;233;234;218mW\033[38;2;238;239;222m&\033[38;2;239;240;223m8\033[38;2;208;209;196ma\033[38;2;188;188;174mp\033[38;2;231;231;215mW\033[38;2;218;218;206m*\033[38;2;144;151;153mQ\033[38;2;109;119;127mz\033[38;2;136;140;144mC\033[38;2;136;142;145mC\033[38;2;62;72;82m1\033[38;2;35;42;59mi\033[38;2;41;45;60mi\033[38;2;41;44;60mi\033[38;2;33;36;47ml\033[38;2;161;142;82mY\033[38;2;190;164;74mC\033[38;2;157;133;51mc\033[38;2;139;116;50mn\033[38;2;138;116;49mn\033[38;2;141;115;50mn\033[38;2;142;118;53mu\033[38;2;150;126;52mv\033[38;2;150;125;51mv\033[38;2;151;125;50mv\033[38;2;146;122;46mu\033[38;2;146;134;95mX\033[38;2;129;132;125mY\033[38;2;32;35;48ml\033[38;2;36;37;53m!\033[38;2;38;39;55m!\033[38;2;33;37;52ml\033[38;2;30;33;48ml\033[38;2;39;43;54mi\033[38;2;73;79;84mt\033[38;2;125;129;129mY\033[38;2;135;139;131mJ\033[38;2;61;64;56m_\033[38;2;48;52;43mi\033[38;2;193;194;188mb\033[38;2;255;255;255m$\033[0m                        \033[0m");
  $display("\033[0m                  \033[38;2;255;255;255m$\033[38;2;252;252;251m@\033[38;2;247;245;232m%%\033[38;2;236;237;219m&\033[38;2;234;237;219m&\033[38;2;234;237;218mW\033[38;2;236;238;220m&\033[38;2;233;232;216mW\033[38;2;183;183;170mq\033[38;2;189;190;176md\033[38;2;225;225;208m#\033[38;2;236;238;220m&\033[38;2;235;238;220m&\033[38;2;234;237;220m&\033[38;2;232;235;218mW\033[38;2;233;234;217mW\033[38;2;232;233;217mW\033[38;2;232;234;216mW\033[38;2;235;238;218m&\033[38;2;236;238;219m&\033[38;2;232;235;215mW\033[38;2;234;236;217mW\033[38;2;239;241;222m8\033[38;2;223;226;212m#\033[38;2;186;189;181md\033[38;2;154;157;154m0\033[38;2;103;108;110mu\033[38;2;35;42;55m!\033[38;2;42;47;62m~\033[38;2;42;44;61mi\033[38;2;32;35;47ml\033[38;2;176;156;90mC\033[38;2;239;211;104mp\033[38;2;227;200;93mw\033[38;2;195;171;81mQ\033[38;2;147;128;85mz\033[38;2;149;143;115mJ\033[38;2;136;136;116mY\033[38;2;145;144;114mU\033[38;2;146;137;95mY\033[38;2;146;132;80mz\033[38;2;134;118;68mu\033[38;2;117;106;61mr\033[38;2;144;148;128mC\033[38;2;108;113;108mv\033[38;2;41;43;53mi\033[38;2;29;33;48ml\033[38;2;31;37;52ml\033[38;2;32;36;50ml\033[38;2;61;67;72m-\033[38;2;72;79;79m1\033[38;2;86;90;91mj\033[38;2;83;87;88mj\033[38;2;90;93;86mj\033[38;2;203;203;197mh\033[38;2;255;255;255m$\033[0m                         \033[0m");
  $display("\033[0m                  \033[38;2;255;255;255m$\033[38;2;250;250;247m@\033[38;2;243;242;224m8\033[38;2;235;237;219m&\033[38;2;235;237;217mW\033[38;2;235;236;217mW\033[38;2;237;237;217m&\033[38;2;233;234;215mW\033[38;2;184;187;170mp\033[38;2;206;207;189mh\033[38;2;231;229;211mM\033[38;2;222;220;202m*\033[38;2;236;236;218m&\033[38;2;235;238;221m&\033[38;2;232;235;218mW\033[38;2;232;233;215mW\033[38;2;233;234;216mWWWWW\033[38;2;234;235;216mW\033[38;2;226;227;209m#\033[38;2;214;214;197mo\033[38;2;228;226;213mM\033[38;2;219;216;205m*\033[38;2;112;113;113mv\033[38;2;31;35;51ml\033[38;2;32;40;56m!\033[38;2;57;60;66m_\033[38;2;107;100;71mr\033[38;2;213;190;96mZ\033[38;2;217;198;104mw\033[38;2;183;175;119mO\033[38;2;201;201;175mb\033[38;2;219;220;205m*\033[38;2;203;203;190mh\033[38;2;192;194;180md\033[38;2;159;164;153mO\033[38;2;143;152;147mL\033[38;2;101;116;123mc\033[38;2;73;97;116mx\033[38;2;68;90;114mr\033[38;2;109;121;121mz\033[38;2;167;169;153mZ\033[38;2;146;145;136mC\033[38;2;110;112;106mv\033[38;2;52;56;63m+\033[38;2;31;36;50ml\033[38;2;50;57;65m+\033[38;2;59;67;70m-\033[38;2;99;105;103mn\033[38;2;121;127;119mX\033[38;2;117;118;108mc\033[38;2;205;204;197mh\033[38;2;255;255;255m$\033[0m                         \033[0m");
  $display("\033[0m                  \033[38;2;255;255;255m$\033[38;2;248;247;241mB\033[38;2;236;238;218m&\033[38;2;235;237;218m&\033[38;2;235;235;215mW\033[38;2;236;235;215mW\033[38;2;237;236;216mW\033[38;2;236;237;217m&\033[38;2;188;192;174mp\033[38;2;211;213;193ma\033[38;2;240;238;219m&\033[38;2;223;220;201m*\033[38;2;187;186;168mp\033[38;2;230;231;215mW\033[38;2;234;235;218mW\033[38;2;232;233;215mWW\033[38;2;233;234;216mWWWWW\033[38;2;232;233;215mW\033[38;2;213;214;195mo\033[38;2;198;197;183mb\033[38;2;166;165;156mZ\033[38;2;122;122;117mz\033[38;2;115;117;114mc\033[38;2;141;144;138mC\033[38;2;199;200;189mk\033[38;2;158;164;138m0\033[38;2;160;176;153mZ\033[38;2;130;163;169m0\033[38;2;116;161;186m0\033[38;2;126;168;191mO\033[38;2;139;174;191mm\033[38;2;145;169;177mZ\033[38;2;168;189;194mp\033[38;2;139;165;173mO\033[38;2;100;134;153mY\033[38;2;82;114;138mv\033[38;2;73;101;122mx\033[38;2;72;100;120mx\033[38;2;80;99;112mx\033[38;2;145;151;140mL\033[38;2;160;163;149m0\033[38;2;159;163;150m0\033[38;2;98;100;97mx\033[38;2;35;35;45ml\033[38;2;137;141;131mJ\033[38;2;123;127;115mz\033[38;2;124;127;117mX\033[38;2;127;130;118mX\033[38;2;136;138;124mU\033[38;2;189;189;176mp\033[38;2;255;255;255m$\033[0m                         \033[0m");
  $display("\033[0m                 \033[38;2;255;255;255m$\033[38;2;253;253;255m$\033[38;2;247;247;235mB\033[38;2;233;236;217mW\033[38;2;235;235;217mW\033[38;2;236;235;217mW\033[38;2;234;235;216mW\033[38;2;234;235;217mW\033[38;2;237;238;220m&\033[38;2;200;201;182mk\033[38;2;215;216;198mo\033[38;2;235;237;217mW\033[38;2;226;228;206m#\033[38;2;168;170;150mZ\033[38;2;180;181;163mw\033[38;2;225;224;206m#\033[38;2;235;235;216mW\033[38;2;233;234;215mWW\033[38;2;233;234;216mW\033[38;2;234;235;216mWW\033[38;2;233;234;215mW\033[38;2;232;233;214mW\033[38;2;234;235;216mW\033[38;2;227;229;210mM\033[38;2;223;225;207m#\033[38;2;225;227;207m#\033[38;2;231;231;212mM\033[38;2;240;241;220m&\033[38;2;238;239;217m&\033[38;2;186;200;196mk\033[38;2;121;162;184m0\033[38;2;123;170;193mZ\033[38;2;126;171;193mZ\033[38;2;124;170;192mZ\033[38;2;123;170;192mO\033[38;2;121;166;190mO\033[38;2;105;147;167mJ\033[38;2;122;162;178m0\033[38;2;124;160;173mQ\033[38;2;126;167;181mO\033[38;2;111;147;167mC\033[38;2;89;120;140mc\033[38;2;73;98;120mx\033[38;2;104;115;119mv\033[38;2;140;143;129mJ\033[38;2;109;113;104mv\033[38;2;95;97;90mr\033[38;2;99;103;95mn\033[38;2;141;148;134mC\033[38;2;149;152;132mL\033[38;2;163;165;145m0\033[38;2;162;165;145m0\033[38;2;158;162;143m0\033[38;2;161;164;145m0\033[38;2;241;241;239m%%\033[38;2;255;255;255m$\033[0m                        \033[0m");
  $display("\033[0m                 \033[38;2;255;255;255m$\033[38;2;252;252;249m@\033[38;2;240;239;223m8\033[38;2;241;241;223m8\033[38;2;237;238;221m&\033[38;2;237;237;221m&&\033[38;2;238;239;221m&\033[38;2;240;241;224m8\033[38;2;221;222;206m#\033[38;2;227;228;213mM\033[38;2;236;238;222m&\033[38;2;232;234;217mW\033[38;2;202;204;187mk\033[38;2;198;198;183mb\033[38;2;208;206;190mh\033[38;2;236;235;220m&\033[38;2;238;237;221m&\033[38;2;236;235;218mW\033[38;2;237;237;222m&\033[38;2;238;239;223m&&\033[38;2;237;237;221m&\033[38;2;236;237;221m&\033[38;2;232;233;216mW\033[38;2;205;206;190mh\033[38;2;201;202;187mk\033[38;2;203;205;189mh\033[38;2;222;223;207m#\033[38;2;238;239;225m8\033[38;2;236;236;219m&\033[38;2;237;234;220m&\033[38;2;192;203;202mh\033[38;2;177;199;205mbb\033[38;2;177;200;204mb\033[38;2;176;198;202mb\033[38;2;177;197;200mb\033[38;2;192;199;194mk\033[38;2;214;215;199mo\033[38;2;211;210;191ma\033[38;2;203;206;187mh\033[38;2;197;204;195mh\033[38;2;188;199;198mk\033[38;2;175;184;189mp\033[38;2;166;170;168mm\033[38;2;208;205;192mh\033[38;2;214;212;201mo\033[38;2;218;215;202mo\033[38;2;221;219;207m*\033[38;2;203;204;198mh\033[38;2;206;206;198ma\033[38;2;209;208;200ma\033[38;2;210;212;204mo\033[38;2;209;210;202mo\033[38;2;203;203;193mh\033[38;2;240;240;237m%%\033[38;2;255;255;255m$\033[0m                        \033[0m");
  $display("\033[0m                  \033[38;2;255;255;255m$$\033[38;2;255;255;251m$\033[38;2;255;255;250m$\033[38;2;255;255;255m$$\033[38;2;255;255;250m$\033[38;2;251;251;251m@\033[38;2;255;255;255m$$$$$$$$$\033[38;2;255;255;250m$\033[38;2;255;255;255m$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$$\033[0m                         \033[0m");
endtask

endmodule



